library verilog;
use verilog.vl_types.all;
entity filt_addr_calc_tb is
end filt_addr_calc_tb;
