module adder32b (a, b, cin, s, cout, vdd, gnd);
	input [31:0] a, [31:0] b, cin, vdd, gnd;
	output [31:0] s, cout;