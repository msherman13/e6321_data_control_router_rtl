module dc_router_top (
	chipselect, 
	clk, 
	reset, 
	instruction, 
	offset, 
	filesize, 
	acc_done, 
	fft_enable, 
	fir_enable, 
	iir_enable, 
	data_bus, 
	fft_data_in, 
	fir_data_in, 
	iir_data_in, 
	fft_data_out, 
	fir_data_out, 
	iir_data_out, 
	to_fft_empty, 
	to_fft_full, 
	from_fft_empty, 
	from_fft_full, 
	to_fir_empty, 
	to_fir_full, 
	from_fir_empty, 
	from_fir_full, 
	to_iir_empty, 
	to_iir_full, 
	from_iir_empty, 
	from_iir_full, 
	fft_put_req, 
	fft_get_req, 
	fir_put_req, 
	fir_get_req, 
	iir_put_req, 
	iir_get_req, 
	ram_read_enable, 
	ram_write_enable, 
	addr);
   input chipselect;
   input clk;
   input reset;
   input [31:0] instruction;
   input [31:0] offset;
   input [31:0] filesize;
   output acc_done;
   output fft_enable;
   output fir_enable;
   output iir_enable;
   inout [31:0] data_bus;
   input [31:0] fft_data_in;
   input [31:0] fir_data_in;
   input [31:0] iir_data_in;
   output [31:0] fft_data_out;
   output [31:0] fir_data_out;
   output [31:0] iir_data_out;
   input to_fft_empty;
   input to_fft_full;
   input from_fft_empty;
   input from_fft_full;
   input to_fir_empty;
   input to_fir_full;
   input from_fir_empty;
   input from_fir_full;
   input to_iir_empty;
   input to_iir_full;
   input from_iir_empty;
   input from_iir_full;
   output fft_put_req;
   output fft_get_req;
   output fir_put_req;
   output fir_get_req;
   output iir_put_req;
   output iir_get_req;
   output ram_read_enable;
   output ram_write_enable;
   output [31:0] addr;

   // Internal wires
   wire clk__L1_N0;
   wire FE_OCP_RBN1982_add_x_19_4_n157;
   wire FE_OCP_RBN1981_add_x_19_4_n157;
   wire FE_OCP_RBN1980_add_x_19_4_n178;
   wire FE_OCP_RBN1979_add_x_19_4_n178;
   wire FE_OCP_RBN1978_add_x_19_4_n178;
   wire FE_OCP_RBN1974_offset_1_;
   wire FE_OCP_RBN1973_offset_1_;
   wire FE_OCP_DRV_N1968_filesize_8_;
   wire FE_RN_468_0;
   wire FE_RN_467_0;
   wire FE_RN_459_0;
   wire FE_RN_458_0;
   wire FE_RN_450_0;
   wire FE_RN_449_0;
   wire FE_RN_448_0;
   wire FE_RN_447_0;
   wire FE_RN_446_0;
   wire FE_RN_445_0;
   wire FE_RN_444_0;
   wire FE_RN_443_0;
   wire FE_RN_438_0;
   wire FE_RN_437_0;
   wire FE_OCP_RBN1957_FE_OFN520_add_x_19_1_n157;
   wire FE_OCP_RBN1956_FE_OFN520_add_x_19_1_n157;
   wire FE_OCP_RBN1955_add_x_19_1_n187;
   wire FE_OCPN1947_n1149;
   wire FE_OCPN1945_offset_2_;
   wire FE_OCPN1944_offset_2_;
   wire FE_RN_431_0;
   wire FE_RN_420_0;
   wire FE_RN_419_0;
   wire FE_RN_418_0;
   wire FE_RN_417_0;
   wire FE_RN_416_0;
   wire FE_RN_415_0;
   wire FE_RN_414_0;
   wire FE_RN_413_0;
   wire FE_RN_412_0;
   wire FE_RN_411_0;
   wire FE_RN_410_0;
   wire FE_RN_409_0;
   wire FE_OCPUNCON1943_FE_OFN407_offset_13_;
   wire FE_OCPUNCON1942_FE_OFN399_offset_15_;
   wire FE_OCPUNCON1941_offset_13_;
   wire FE_OCPUNCON1940_offset_15_;
   wire FE_RN_371_0;
   wire FE_OCP_RBN1925_add_x_19_4_n157;
   wire FE_OCP_RBN1919_offset_1_;
   wire FE_OCPN1911_FE_OFN17_n2797;
   wire FE_OCPN1910_n1736;
   wire FE_OCPN1908_add_x_19_3_n136;
   wire FE_OCPN1907_add_x_19_5_n187;
   wire FE_OCPN1906_add_x_19_3_n139;
   wire FE_OCPN1905_FE_OCPUNCON1873_offset_11_;
   wire FE_OCPN1904_FE_OCPUNCON1066_offset_3_;
   wire FE_OCP_DRV_N1894_filesize_29_;
   wire FE_OCPUNCON1888_n2813;
   wire FE_OCPUNCON1887_n2813;
   wire FE_OCPUNCON1886_n2813;
   wire FE_OCPUNCON1885_n2813;
   wire FE_OCPUNCON1884_n2813;
   wire FE_OCPUNCON1883_n2813;
   wire FE_OCPUNCON1882_n2813;
   wire FE_OCPUNCON1881_n2813;
   wire FE_OCPUNCON1880_n2787;
   wire FE_OCPUNCON1879_n2813;
   wire FE_OCPUNCON1878_n2787;
   wire FE_OCPUNCON1877_FE_OFN374_offset_22_;
   wire FE_OCPUNCON1876_offset_22_;
   wire FE_OCPUNCON1875_offset_4_;
   wire FE_OCPUNCON1874_offset_1_;
   wire FE_OCPUNCON1873_offset_11_;
   wire FE_RN_368_0;
   wire FE_RN_367_0;
   wire FE_OCP_DRV_N1872_filesize_18_;
   wire FE_RN_349_0;
   wire FE_RN_348_0;
   wire FE_RN_347_0;
   wire FE_RN_346_0;
   wire FE_RN_345_0;
   wire FE_RN_344_0;
   wire FE_RN_343_0;
   wire FE_RN_342_0;
   wire FE_RN_341_0;
   wire FE_RN_340_0;
   wire FE_RN_339_0;
   wire FE_RN_338_0;
   wire FE_OCP_RBN1842_offset_7_;
   wire FE_OCP_RBN1841_offset_7_;
   wire FE_OCP_RBN1840_offset_7_;
   wire FE_OCPN1825_add_x_19_3_n68;
   wire FE_OCP_DRV_N1824_filesize_19_;
   wire FE_OCP_DRV_N1818_filesize_20_;
   wire FE_RN_310_0;
   wire FE_OCP_RBN1788_add_x_19_3_n163;
   wire FE_OCP_RBN1787_add_x_19_3_n163;
   wire FE_OCPUNCON1750_offset_1_;
   wire FE_OCPN1732_n1718;
   wire FE_OCPN1731_FE_OCPUNCON1650_add_x_19_4_n43;
   wire FE_OCPN1730_add_x_19_0_n43;
   wire FE_OCPN1729_FE_OFN528_add_x_19_0_n113;
   wire FE_OCPN1728_FE_OFN528_add_x_19_0_n113;
   wire FE_OCPUNCON1686_offset_20_;
   wire FE_OCPUNCON1684_offset_6_;
   wire FE_RN_304_0;
   wire FE_RN_303_0;
   wire FE_RN_302_0;
   wire FE_RN_301_0;
   wire FE_RN_294_0;
   wire FE_RN_293_0;
   wire FE_RN_292_0;
   wire FE_RN_291_0;
   wire FE_RN_290_0;
   wire FE_RN_289_0;
   wire FE_RN_285_0;
   wire FE_RN_284_0;
   wire FE_RN_269_0;
   wire FE_RN_241_0;
   wire FE_RN_240_0;
   wire FE_RN_239_0;
   wire FE_RN_238_0;
   wire FE_RN_237_0;
   wire FE_RN_219_0;
   wire FE_RN_218_0;
   wire FE_RN_217_0;
   wire FE_RN_214_0;
   wire FE_RN_213_0;
   wire FE_OCPUNCON1650_add_x_19_4_n43;
   wire FE_RN_212_0;
   wire FE_RN_208_0;
   wire FE_RN_207_0;
   wire FE_OCPUNCON1576_n2812;
   wire FE_OCPUNCON1575_n2812;
   wire FE_OCPUNCON1574_n2812;
   wire FE_OCPUNCON1573_n2812;
   wire FE_OCPUNCON1572_n2812;
   wire FE_OCPUNCON1571_n2812;
   wire FE_OCPUNCON1570_n2812;
   wire FE_OCPUNCON1569_n2812;
   wire FE_OCPUNCON1568_n2812;
   wire FE_OCPUNCON1567_n1717;
   wire FE_OCPUNCON1566_n1789;
   wire FE_OCPUNCON1565_n1789;
   wire FE_OCPUNCON1564_offset_5_;
   wire FE_OCPUNCON1563_offset_3_;
   wire FE_OCPUNCON1562_filesize_10_;
   wire FE_RN_205_0;
   wire FE_RN_203_0;
   wire FE_RN_202_0;
   wire FE_RN_201_0;
   wire FE_RN_200_0;
   wire FE_RN_199_0;
   wire FE_RN_198_0;
   wire FE_RN_197_0;
   wire FE_RN_192_0;
   wire FE_RN_191_0;
   wire FE_RN_190_0;
   wire FE_RN_188_0;
   wire FE_RN_187_0;
   wire FE_OCP_RBN1495_offset_5_;
   wire FE_OCP_RBN1494_offset_5_;
   wire FE_OCP_RBN1493_offset_5_;
   wire FE_OCP_RBN1492_offset_5_;
   wire FE_OCPUNCON1425_FE_OFN443_offset_4_;
   wire FE_OCP_DRV_N1389_filesize_16_;
   wire FE_OCP_RBN1383_add_x_19_0_n92;
   wire FE_OCP_RBN1381_add_x_19_3_n92;
   wire FE_OCP_RBN1379_add_x_19_1_n69;
   wire FE_OCP_RBN1378_add_x_19_3_n113;
   wire FE_OCP_RBN1366_FE_OCP_DRV_N1167_offset_20_;
   wire FE_OCP_RBN1365_FE_OCP_DRV_N1167_offset_20_;
   wire FE_OCP_RBN1364_FE_OCP_DRV_N1167_offset_20_;
   wire FE_OCP_RBN1363_FE_OCP_DRV_N1167_offset_20_;
   wire FE_OCPN1362_add_x_19_2_n83;
   wire FE_OCP_DRV_N1336_filesize_0_;
   wire FE_OCPUNCON1318_FE_OFN361_offset_25_;
   wire FE_OCPUNCON1278_offset_7_;
   wire FE_OCPN1257_add_x_19_0_n162;
   wire FE_OCPN1256_add_x_19_3_n162;
   wire FE_OCPN1255_add_x_19_3_n181;
   wire FE_OCPN1230_n1611;
   wire FE_OCPN1229_add_x_19_5_n68;
   wire FE_OCPN1226_add_x_19_4_n112;
   wire FE_OCPN1225_add_x_19_5_n170;
   wire FE_OCPN1224_FE_OFN445_offset_4_;
   wire FE_OCPN1223_add_x_19_1_n181;
   wire FE_OCPN1222_add_x_19_5_n162;
   wire FE_OCPN1221_add_x_19_4_n162;
   wire FE_OCPN1220_add_x_19_2_n181;
   wire FE_OCPN1189_add_x_19_0_n181;
   wire FE_OCPN1188_offset_3_;
   wire FE_OCP_DRV_N1099_filesize_14_;
   wire FE_OCPUNCON1093_n2805;
   wire FE_OCPUNCON1092_n2805;
   wire FE_OCPUNCON1091_n2805;
   wire FE_OCPUNCON1090_n2805;
   wire FE_OCPUNCON1089_n2805;
   wire FE_OCPUNCON1088_n2805;
   wire FE_OCPUNCON1087_n2805;
   wire FE_OCPUNCON1086_n2805;
   wire FE_OCPUNCON1085_n2805;
   wire FE_OCPUNCON1084_n2805;
   wire FE_OCPUNCON1083_n2805;
   wire FE_OCPUNCON1082_n2589;
   wire FE_OCPUNCON1081_n2589;
   wire FE_OCPUNCON1080_FE_OFN386_offset_18_;
   wire FE_OCPUNCON1079_FE_OFN382_offset_19_;
   wire FE_OCPUNCON1078_FE_OFN377_offset_21_;
   wire FE_OCPUNCON1077_FE_OFN459_offset_0_;
   wire FE_OCPUNCON1076_FE_OFN451_offset_2_;
   wire FE_OCPUNCON1075_FE_OFN447_offset_3_;
   wire FE_OCPUNCON1073_FE_OFN410_offset_12_;
   wire FE_OCPUNCON1072_FE_OFN386_offset_18_;
   wire FE_OCPUNCON1071_FE_OFN382_offset_19_;
   wire FE_OCPUNCON1070_FE_OFN377_offset_21_;
   wire FE_OCPUNCON1069_FE_OFN369_offset_23_;
   wire FE_OCPUNCON1068_offset_0_;
   wire FE_OCPUNCON1066_offset_3_;
   wire FE_OCPUNCON1065_offset_2_;
   wire FE_OCPUNCON1062_offset_19_;
   wire FE_OCPUNCON1060_offset_21_;
   wire FE_OCPUNCON1058_filesize_3_;
   wire FE_RN_184_0;
   wire FE_RN_183_0;
   wire FE_RN_182_0;
   wire FE_RN_181_0;
   wire FE_RN_176_0;
   wire FE_RN_175_0;
   wire FE_RN_174_0;
   wire FE_RN_173_0;
   wire FE_RN_168_0;
   wire FE_RN_167_0;
   wire FE_RN_166_0;
   wire FE_RN_165_0;
   wire FE_RN_164_0;
   wire FE_RN_163_0;
   wire FE_RN_162_0;
   wire FE_RN_161_0;
   wire FE_RN_158_0;
   wire FE_RN_157_0;
   wire FE_RN_156_0;
   wire FE_RN_155_0;
   wire FE_RN_154_0;
   wire FE_RN_153_0;
   wire FE_RN_152_0;
   wire FE_RN_149_0;
   wire FE_RN_146_0;
   wire FE_RN_145_0;
   wire FE_RN_144_0;
   wire FE_RN_143_0;
   wire FE_RN_142_0;
   wire FE_RN_136_0;
   wire FE_RN_135_0;
   wire FE_RN_134_0;
   wire FE_RN_132_0;
   wire FE_RN_129_0;
   wire FE_RN_128_0;
   wire FE_RN_113_0;
   wire FE_RN_112_0;
   wire FE_RN_111_0;
   wire FE_RN_110_0;
   wire FE_RN_109_0;
   wire FE_RN_108_0;
   wire FE_RN_107_0;
   wire FE_RN_106_0;
   wire FE_RN_105_0;
   wire FE_RN_104_0;
   wire FE_RN_103_0;
   wire FE_RN_102_0;
   wire FE_RN_101_0;
   wire FE_RN_100_0;
   wire FE_RN_99_0;
   wire FE_RN_98_0;
   wire FE_RN_92_0;
   wire FE_RN_91_0;
   wire FE_RN_87_0;
   wire FE_RN_86_0;
   wire FE_RN_85_0;
   wire FE_RN_84_0;
   wire FE_RN_64_0;
   wire FE_RN_59_0;
   wire FE_RN_56_0;
   wire FE_RN_55_0;
   wire FE_RN_46_0;
   wire FE_RN_45_0;
   wire FE_RN_41_0;
   wire FE_RN_40_0;
   wire FE_RN_39_0;
   wire FE_RN_38_0;
   wire FE_RN_35_0;
   wire FE_RN_34_0;
   wire FE_RN_33_0;
   wire FE_RN_32_0;
   wire FE_RN_31_0;
   wire FE_RN_30_0;
   wire FE_RN_29_0;
   wire FE_RN_28_0;
   wire FE_RN_7_0;
   wire FE_RN_6_0;
   wire FE_RN_5_0;
   wire FE_RN_2_0;
   wire FE_RN_1_0;
   wire FE_RN_0_0;
   wire FE_OCPUNCON726_FE_OFN435_offset_6_;
   wire FE_OCPUNCON658_FE_OFN422_offset_9_;
   wire FE_OCPUNCON657_FE_OFN418_offset_10_;
   wire FE_OCPUNCON656_FE_OFN414_offset_11_;
   wire FE_OCPUNCON654_FE_OFN422_offset_9_;
   wire FE_OCPUNCON653_FE_OFN418_offset_10_;
   wire FE_OCPUNCON652_FE_OFN414_offset_11_;
   wire FE_OFN615_filesize_0_;
   wire FE_OFN614_filesize_1_;
   wire FE_OFN613_filesize_2_;
   wire FE_OFN612_filesize_4_;
   wire FE_OFN611_filesize_5_;
   wire FE_OFN610_filesize_6_;
   wire FE_OFN609_filesize_7_;
   wire FE_OFN608_filesize_8_;
   wire FE_OFN607_filesize_9_;
   wire FE_OFN605_filesize_11_;
   wire FE_OFN604_filesize_12_;
   wire FE_OFN603_filesize_13_;
   wire FE_OFN602_filesize_14_;
   wire FE_OFN600_filesize_17_;
   wire FE_OFN599_filesize_18_;
   wire FE_OFN598_filesize_19_;
   wire FE_OFN597_filesize_20_;
   wire FE_OFN596_filesize_21_;
   wire FE_OFN595_filesize_24_;
   wire FE_OFN594_filesize_26_;
   wire FE_OFN593_filesize_27_;
   wire FE_OFN592_filesize_28_;
   wire FE_OFN591_filesize_29_;
   wire FE_OFN580_offset_16_;
   wire FE_OFN568_offset_28_;
   wire FE_OFN567_n2070;
   wire FE_OFN566_n2066;
   wire FE_OFN565_n2066;
   wire FE_OFN564_n2066;
   wire FE_OFN563_n2060;
   wire FE_OFN562_n2060;
   wire FE_OFN561_n2587;
   wire FE_OFN560_n2587;
   wire FE_OFN559_offset_30_;
   wire FE_OFN558_n2441;
   wire FE_OFN557_n2441;
   wire FE_OFN553_n1789;
   wire FE_OFN552_n1751;
   wire FE_OFN551_n1751;
   wire FE_OFN550_n1750;
   wire FE_OFN549_n1763;
   wire FE_OFN548_n1763;
   wire FE_OFN547_n2803;
   wire FE_OFN545_addr_calc_iir_write_addr_11_;
   wire FE_OFN544_addr_calc_fft_read_addr_11_;
   wire FE_OFN543_addr_calc_fir_write_addr_17_;
   wire FE_OFN541_addr_calc_iir_read_addr_9_;
   wire FE_OFN540_DP_OP_158_296_6262_n765;
   wire FE_OFN539_DP_OP_158_296_6262_n318;
   wire FE_OFN538_DP_OP_158_296_6262_n1659;
   wire FE_OFN537_DP_OP_159_297_3515_n301;
   wire FE_OFN536_addr_calc_iir_read_addr_7_;
   wire FE_OFN535_DP_OP_159_297_3515_n726;
   wire FE_OFN534_addr_calc_iir_write_addr_7_;
   wire FE_OFN533_addr_calc_fir_write_addr_7_;
   wire FE_OFN532_addr_calc_fft_read_addr_7_;
   wire FE_OFN531_add_x_19_5_n43;
   wire FE_OFN529_DP_OP_158_296_6262_n838;
   wire FE_OFN528_add_x_19_0_n113;
   wire FE_OFN527_add_x_19_4_n113;
   wire FE_OFN526_add_x_19_2_n113;
   wire FE_OFN525_add_x_19_3_n157;
   wire FE_OFN524_n1659;
   wire FE_OFN523_add_x_19_1_n113;
   wire FE_OFN522_add_x_19_5_n114;
   wire FE_OFN521_n1592;
   wire FE_OFN520_add_x_19_1_n157;
   wire FE_OFN519_DP_OP_159_297_3515_n1039;
   wire FE_OFN518_n2372;
   wire FE_OFN517_addr_calc_fft_read_calc_count_0_;
   wire FE_OFN516_from_iir_full;
   wire FE_OFN515_from_iir_empty;
   wire FE_OFN514_to_iir_full;
   wire FE_OFN513_to_iir_empty;
   wire FE_OFN512_from_fir_full;
   wire FE_OFN511_from_fir_empty;
   wire FE_OFN510_to_fir_full;
   wire FE_OFN509_to_fir_empty;
   wire FE_OFN508_from_fft_full;
   wire FE_OFN507_from_fft_empty;
   wire FE_OFN506_to_fft_full;
   wire FE_OFN505_to_fft_empty;
   wire FE_OFN504_iir_data_in_9_;
   wire FE_OFN503_fft_data_in_9_;
   wire FE_OFN502_filesize_0_;
   wire FE_OFN501_filesize_1_;
   wire FE_OFN500_filesize_1_;
   wire FE_OFN499_filesize_2_;
   wire FE_OFN498_filesize_3_;
   wire FE_OFN496_filesize_4_;
   wire FE_OFN495_filesize_5_;
   wire FE_OFN494_filesize_6_;
   wire FE_OFN493_filesize_7_;
   wire FE_OFN492_filesize_8_;
   wire FE_OFN491_filesize_9_;
   wire FE_OFN490_filesize_10_;
   wire FE_OFN489_filesize_11_;
   wire FE_OFN488_filesize_12_;
   wire FE_OFN487_filesize_13_;
   wire FE_OFN486_filesize_14_;
   wire FE_OFN485_filesize_14_;
   wire FE_OFN484_filesize_15_;
   wire FE_OFN483_filesize_15_;
   wire FE_OFN482_filesize_16_;
   wire FE_OFN481_filesize_16_;
   wire FE_OFN480_filesize_17_;
   wire FE_OFN479_filesize_18_;
   wire FE_OFN478_filesize_19_;
   wire FE_OFN477_filesize_20_;
   wire FE_OFN476_filesize_21_;
   wire FE_OFN475_filesize_22_;
   wire FE_OFN474_filesize_22_;
   wire FE_OFN473_filesize_23_;
   wire FE_OFN472_filesize_23_;
   wire FE_OFN471_filesize_24_;
   wire FE_OFN470_filesize_25_;
   wire FE_OFN469_filesize_25_;
   wire FE_OFN468_filesize_26_;
   wire FE_OFN467_filesize_27_;
   wire FE_OFN466_filesize_28_;
   wire FE_OFN465_filesize_29_;
   wire FE_OFN464_filesize_29_;
   wire FE_OFN463_filesize_30_;
   wire FE_OFN462_filesize_31_;
   wire FE_OFN461_offset_0_;
   wire FE_OFN459_offset_0_;
   wire FE_OFN452_offset_2_;
   wire FE_OFN451_offset_2_;
   wire FE_OFN449_offset_3_;
   wire FE_OFN447_offset_3_;
   wire FE_OFN444_offset_4_;
   wire FE_OFN443_offset_4_;
   wire FE_OFN436_offset_6_;
   wire FE_OFN435_offset_6_;
   wire FE_OFN429_offset_8_;
   wire FE_OFN428_offset_8_;
   wire FE_OFN427_offset_8_;
   wire FE_OFN426_offset_8_;
   wire FE_OFN424_offset_9_;
   wire FE_OFN422_offset_9_;
   wire FE_OFN421_offset_10_;
   wire FE_OFN418_offset_10_;
   wire FE_OFN417_offset_11_;
   wire FE_OFN413_offset_12_;
   wire FE_OFN411_offset_12_;
   wire FE_OFN410_offset_12_;
   wire FE_OFN408_offset_13_;
   wire FE_OFN407_offset_13_;
   wire FE_OFN405_offset_14_;
   wire FE_OFN404_offset_14_;
   wire FE_OFN403_offset_14_;
   wire FE_OFN402_offset_14_;
   wire FE_OFN400_offset_15_;
   wire FE_OFN399_offset_15_;
   wire FE_OFN397_offset_16_;
   wire FE_OFN396_offset_16_;
   wire FE_OFN395_offset_16_;
   wire FE_OFN394_offset_16_;
   wire FE_OFN393_offset_17_;
   wire FE_OFN392_offset_17_;
   wire FE_OFN391_offset_17_;
   wire FE_OFN390_offset_17_;
   wire FE_OFN389_offset_18_;
   wire FE_OFN386_offset_18_;
   wire FE_OFN384_offset_19_;
   wire FE_OFN382_offset_19_;
   wire FE_OFN380_offset_21_;
   wire FE_OFN377_offset_21_;
   wire FE_OFN375_offset_22_;
   wire FE_OFN374_offset_22_;
   wire FE_OFN372_offset_23_;
   wire FE_OFN371_offset_23_;
   wire FE_OFN369_offset_23_;
   wire FE_OFN368_offset_24_;
   wire FE_OFN367_offset_24_;
   wire FE_OFN366_offset_24_;
   wire FE_OFN365_offset_24_;
   wire FE_OFN364_offset_25_;
   wire FE_OFN363_offset_25_;
   wire FE_OFN361_offset_25_;
   wire FE_OFN360_offset_26_;
   wire FE_OFN359_offset_26_;
   wire FE_OFN358_offset_26_;
   wire FE_OFN357_offset_26_;
   wire FE_OFN356_offset_27_;
   wire FE_OFN355_offset_27_;
   wire FE_OFN354_offset_27_;
   wire FE_OFN353_offset_27_;
   wire FE_OFN352_offset_28_;
   wire FE_OFN351_offset_28_;
   wire FE_OFN350_offset_28_;
   wire FE_OFN349_offset_28_;
   wire FE_OFN348_offset_29_;
   wire FE_OFN347_offset_29_;
   wire FE_OFN346_offset_29_;
   wire FE_OFN345_offset_29_;
   wire FE_OFN344_offset_30_;
   wire FE_OFN343_offset_30_;
   wire FE_OFN341_offset_30_;
   wire FE_OFN340_offset_31_;
   wire FE_OFN339_offset_31_;
   wire FE_OFN338_offset_31_;
   wire FE_OFN337_offset_31_;
   wire FE_OFN336_instruction_0_;
   wire FE_OFN335_instruction_2_;
   wire FE_OFN334_data_to_fft;
   wire FE_OFN333_data_to_fft;
   wire FE_OFN332_data_cntl_N63;
   wire FE_OFN331_data_to_fir;
   wire FE_OFN330_data_to_fir;
   wire FE_OFN329_data_cntl_N99;
   wire FE_OFN328_data_to_iir;
   wire FE_OFN327_data_to_iir;
   wire FE_OFN326_data_cntl_N191;
   wire FE_OFN325_data_from_fft;
   wire FE_OFN324_data_from_fft;
   wire FE_OFN323_data_from_fft;
   wire FE_OFN322_data_cntl_N9;
   wire FE_OFN321_data_from_fir;
   wire FE_OFN320_data_from_fir;
   wire FE_OFN319_data_from_fir;
   wire FE_OFN318_data_cntl_N95;
   wire FE_OFN317_data_from_iir;
   wire FE_OFN316_data_from_iir;
   wire FE_OFN315_data_from_iir;
   wire FE_OFN314_data_cntl_N159;
   wire FE_OFN313_n2643;
   wire FE_OFN312_n2643;
   wire FE_OFN311_n2643;
   wire FE_OFN310_n2643;
   wire FE_OFN309_n2644;
   wire FE_OFN308_n2644;
   wire FE_OFN307_n2644;
   wire FE_OFN306_n2644;
   wire FE_OFN305_n2645;
   wire FE_OFN304_n2645;
   wire FE_OFN303_n2645;
   wire FE_OFN302_n2645;
   wire FE_OFN301_n2646;
   wire FE_OFN300_n2646;
   wire FE_OFN299_n2646;
   wire FE_OFN298_n2646;
   wire FE_OFN297_n2642;
   wire FE_OFN296_n2642;
   wire FE_OFN295_n2642;
   wire FE_OFN294_n2642;
   wire FE_OFN293_n2641;
   wire FE_OFN292_n2641;
   wire FE_OFN291_n2641;
   wire FE_OFN290_n2641;
   wire FE_OFN289_n2641;
   wire FE_OFN288_addr_calc_fft_read_calc_count_21_;
   wire FE_OFN287_addr_calc_fft_read_calc_count_17_;
   wire FE_OFN286_addr_calc_iir_read_calc_count_30_;
   wire FE_OFN285_addr_calc_fft_write_calc_count_22_;
   wire FE_OFN284_addr_calc_fft_write_calc_count_22_;
   wire FE_OFN283_addr_calc_fir_write_calc_count_20_;
   wire FE_OFN282_addr_calc_fir_write_calc_count_20_;
   wire FE_OFN281_addr_calc_fft_write_calc_count_20_;
   wire FE_OFN280_addr_calc_fft_write_calc_count_20_;
   wire FE_OFN279_addr_calc_fft_write_calc_count_30_;
   wire FE_OFN278_addr_calc_fft_read_calc_count_30_;
   wire FE_OFN277_addr_calc_fft_write_calc_count_24_;
   wire FE_OFN276_addr_calc_fft_write_calc_count_24_;
   wire FE_OFN275_addr_calc_fft_read_calc_count_29_;
   wire FE_OFN274_addr_calc_fft_write_calc_count_31_;
   wire FE_OFN273_addr_calc_fir_write_calc_count_29_;
   wire FE_OFN272_addr_calc_fft_write_calc_count_6_;
   wire FE_OFN271_addr_calc_fft_write_calc_count_6_;
   wire FE_OFN270_addr_calc_fir_read_calc_count_26_;
   wire FE_OFN269_addr_calc_fir_read_calc_count_26_;
   wire FE_OFN268_addr_calc_fir_write_calc_count_26_;
   wire FE_OFN267_addr_calc_fir_write_calc_count_26_;
   wire FE_OFN266_addr_calc_iir_write_calc_count_18_;
   wire FE_OFN265_addr_calc_iir_write_calc_count_18_;
   wire FE_OFN264_addr_calc_fft_read_calc_count_4_;
   wire FE_OFN263_addr_calc_fft_read_calc_count_4_;
   wire FE_OFN262_addr_calc_fir_write_calc_count_31_;
   wire FE_OFN261_addr_calc_fir_read_calc_count_31_;
   wire FE_OFN260_addr_calc_fft_write_calc_count_0_;
   wire FE_OFN259_addr_calc_fft_write_calc_count_14_;
   wire FE_OFN258_addr_calc_fft_write_calc_count_14_;
   wire FE_OFN257_addr_calc_fir_write_calc_count_8_;
   wire FE_OFN256_addr_calc_fir_write_calc_count_8_;
   wire FE_OFN255_addr_calc_fir_write_calc_count_8_;
   wire FE_OFN254_addr_calc_fir_write_calc_count_6_;
   wire FE_OFN253_addr_calc_fir_write_calc_count_6_;
   wire FE_OFN252_addr_calc_fir_write_calc_count_0_;
   wire FE_OFN251_addr_calc_fft_read_calc_count_5_;
   wire FE_OFN250_addr_calc_iir_write_calc_count_3_;
   wire FE_OFN249_addr_calc_fir_read_calc_count_1_;
   wire FE_OFN248_addr_calc_iir_read_calc_count_10_;
   wire FE_OFN247_addr_calc_iir_read_calc_count_7_;
   wire FE_OFN246_addr_calc_iir_read_calc_count_7_;
   wire FE_OFN245_addr_calc_fir_read_calc_count_5_;
   wire FE_OFN244_addr_calc_iir_read_calc_count_4_;
   wire FE_OFN243_addr_calc_fir_read_calc_count_27_;
   wire FE_OFN242_addr_calc_fir_write_calc_count_1_;
   wire FE_OFN241_addr_calc_fir_write_calc_count_4_;
   wire FE_OFN240_addr_calc_iir_write_calc_count_31_;
   wire FE_OFN239_addr_calc_iir_write_calc_count_30_;
   wire FE_OFN238_addr_calc_fir_write_calc_count_30_;
   wire FE_OFN237_addr_calc_iir_read_calc_count_11_;
   wire FE_OFN236_addr_calc_iir_read_calc_count_11_;
   wire FE_OFN235_addr_calc_iir_read_calc_count_27_;
   wire FE_OFN234_addr_calc_iir_read_calc_count_31_;
   wire FE_OFN233_addr_calc_fir_write_calc_count_12_;
   wire FE_OFN232_addr_calc_fir_write_calc_count_12_;
   wire FE_OFN231_addr_calc_fir_write_calc_count_25_;
   wire FE_OFN230_addr_calc_iir_write_calc_count_15_;
   wire FE_OFN229_addr_calc_iir_write_calc_count_15_;
   wire FE_OFN228_fft_enable;
   wire FE_OFN227_addr_calc_fir_read_calc_count_7_;
   wire FE_OFN226_addr_calc_fft_read_calc_count_31_;
   wire FE_OFN225_addr_calc_fft_read_calc_count_6_;
   wire FE_OFN224_addr_calc_fft_read_calc_count_6_;
   wire FE_OFN223_n643;
   wire FE_OFN222_n643;
   wire FE_OFN221_n643;
   wire FE_OFN220_n643;
   wire FE_OFN219_n643;
   wire FE_OFN218_n643;
   wire FE_OFN217_n643;
   wire FE_OFN216_n643;
   wire FE_OFN215_n643;
   wire FE_OFN214_n515;
   wire FE_OFN213_n515;
   wire FE_OFN212_n515;
   wire FE_OFN211_n515;
   wire FE_OFN210_n515;
   wire FE_OFN209_n515;
   wire FE_OFN208_n515;
   wire FE_OFN207_n515;
   wire FE_OFN206_n387;
   wire FE_OFN205_n387;
   wire FE_OFN204_n387;
   wire FE_OFN203_n387;
   wire FE_OFN202_n387;
   wire FE_OFN201_n387;
   wire FE_OFN200_n387;
   wire FE_OFN199_n387;
   wire FE_OFN198_n387;
   wire FE_OFN197_n387;
   wire FE_OFN196_n707;
   wire FE_OFN195_n707;
   wire FE_OFN194_n707;
   wire FE_OFN193_n707;
   wire FE_OFN192_n707;
   wire FE_OFN191_n707;
   wire FE_OFN190_n707;
   wire FE_OFN189_n579;
   wire FE_OFN188_n579;
   wire FE_OFN187_n579;
   wire FE_OFN186_n579;
   wire FE_OFN185_n579;
   wire FE_OFN184_n579;
   wire FE_OFN183_n579;
   wire FE_OFN182_n451;
   wire FE_OFN181_n451;
   wire FE_OFN180_n451;
   wire FE_OFN179_n451;
   wire FE_OFN178_n451;
   wire FE_OFN177_n451;
   wire FE_OFN176_n451;
   wire FE_OFN175_n131;
   wire FE_OFN174_n131;
   wire FE_OFN173_n131;
   wire FE_OFN172_n131;
   wire FE_OFN171_n195;
   wire FE_OFN170_n195;
   wire FE_OFN169_n195;
   wire FE_OFN168_n195;
   wire FE_OFN167_n259;
   wire FE_OFN166_n259;
   wire FE_OFN165_n259;
   wire FE_OFN164_n259;
   wire FE_OFN163_n323;
   wire FE_OFN162_n323;
   wire FE_OFN161_n323;
   wire FE_OFN160_n323;
   wire FE_OFN159_n67;
   wire FE_OFN158_n67;
   wire FE_OFN157_n67;
   wire FE_OFN156_n67;
   wire FE_OFN155_n3;
   wire FE_OFN154_n3;
   wire FE_OFN153_n3;
   wire FE_OFN152_n3;
   wire FE_OFN151_n2074;
   wire FE_OFN150_add_x_22_4_n59;
   wire FE_OFN149_add_x_22_5_n94;
   wire FE_OFN148_add_x_22_5_n59;
   wire FE_OFN147_add_x_22_2_n59;
   wire FE_OFN146_n801;
   wire FE_OFN145_n801;
   wire FE_OFN144_add_x_19_5_n59;
   wire FE_OFN143_add_x_19_3_n59;
   wire FE_OFN142_add_x_19_2_n59;
   wire FE_OFN140_add_x_19_5_n115;
   wire FE_OFN139_add_x_19_0_n157;
   wire FE_OFN137_addr_calc_fft_read_addr_10_;
   wire FE_OFN136_addr_calc_fft_read_addr_29_;
   wire FE_OFN135_addr_calc_fft_read_addr_30_;
   wire FE_OFN133_addr_calc_fft_read_addr_28_;
   wire FE_OFN132_addr_calc_fir_write_addr_4_;
   wire FE_OFN131_addr_calc_fir_write_addr_16_;
   wire FE_OFN129_add_x_19_5_n157;
   wire FE_OFN128_addr_calc_iir_write_addr_10_;
   wire FE_OFN127_addr_calc_iir_write_addr_9_;
   wire FE_OFN126_addr_calc_iir_write_addr_25_;
   wire FE_OFN125_addr_calc_iir_write_addr_19_;
   wire FE_OFN124_addr_calc_iir_write_addr_16_;
   wire FE_OFN123_addr_calc_iir_write_addr_21_;
   wire FE_OFN122_add_x_19_2_n157;
   wire FE_OFN121_addr_calc_iir_read_addr_4_;
   wire FE_OFN118_addr_calc_iir_read_addr_15_;
   wire FE_OFN117_addr_calc_iir_read_addr_10_;
   wire FE_OFN116_addr_calc_iir_read_addr_24_;
   wire FE_OFN114_DP_OP_159_297_3515_n852;
   wire FE_OFN113_DP_OP_158_296_6262_n1791;
   wire FE_OFN112_DP_OP_158_296_6262_n1791;
   wire FE_OFN93_n1192;
   wire FE_OFN92_n1192;
   wire FE_OFN91_n1192;
   wire FE_OFN90_n1192;
   wire FE_OFN89_n2654;
   wire FE_OFN88_n2654;
   wire FE_OFN87_n2654;
   wire FE_OFN86_n2654;
   wire FE_OFN85_n2654;
   wire FE_OFN84_n2787;
   wire FE_OFN83_n2787;
   wire FE_OFN82_n2787;
   wire FE_OFN81_n2787;
   wire FE_OFN80_n2787;
   wire FE_OFN79_n2787;
   wire FE_OFN78_n2787;
   wire FE_OFN75_n2599;
   wire FE_OFN71_n2809;
   wire FE_OFN70_n2809;
   wire FE_OFN69_n2809;
   wire FE_OFN68_n2809;
   wire FE_OFN67_n2809;
   wire FE_OFN66_n2809;
   wire FE_OFN65_n2809;
   wire FE_OFN64_n2809;
   wire FE_OFN63_n2809;
   wire FE_OFN62_n2809;
   wire FE_OFN61_n2807;
   wire FE_OFN60_n2807;
   wire FE_OFN59_n2807;
   wire FE_OFN58_n2807;
   wire FE_OFN57_n2807;
   wire FE_OFN56_n2807;
   wire FE_OFN55_n2807;
   wire FE_OFN54_n2807;
   wire FE_OFN53_n2807;
   wire FE_OFN52_n2807;
   wire FE_OFN51_n2803;
   wire FE_OFN50_n2803;
   wire FE_OFN49_n2803;
   wire FE_OFN48_n2803;
   wire FE_OFN47_n1758;
   wire FE_OFN35_n2795;
   wire FE_OFN34_n2795;
   wire FE_OFN33_n2795;
   wire FE_OFN32_n2795;
   wire FE_OFN31_n2795;
   wire FE_OFN30_n2795;
   wire FE_OFN29_n2795;
   wire FE_OFN28_n2795;
   wire FE_OFN27_n2795;
   wire FE_OFN26_n2797;
   wire FE_OFN25_n2797;
   wire FE_OFN24_n2797;
   wire FE_OFN23_n2797;
   wire FE_OFN22_n2797;
   wire FE_OFN21_n2797;
   wire FE_OFN20_n2797;
   wire FE_OFN19_n2797;
   wire FE_OFN18_n2797;
   wire FE_OFN17_n2797;
   wire FE_OFN16_n2794;
   wire FE_OFN15_n2794;
   wire FE_OFN14_n2794;
   wire FE_OFN13_n2794;
   wire FE_OFN12_n2794;
   wire FE_OFN11_n2794;
   wire FE_OFN10_n2794;
   wire FE_OFN9_n2794;
   wire FE_OFN8_n2794;
   wire FE_OFN7_n2794;
   wire FE_OFN6_n1750;
   wire FE_OFN4_n1755;
   wire FE_OFN3_n1754;
   wire FE_OFN2_n1754;
   wire FE_OFN1_n1751;
   wire n2814;
   wire n2815;
   wire data_to_fft;
   wire data_from_fft;
   wire data_to_fir;
   wire data_from_fir;
   wire data_to_iir;
   wire data_from_iir;
   wire fft_read_done;
   wire fir_read_done;
   wire fir_write_done;
   wire iir_read_done;
   wire iir_write_done;
   wire fft_put_req_reg;
   wire fir_put_req_reg;
   wire fir_get_req_reg;
   wire iir_put_req_reg;
   wire iir_get_req_reg;
   wire \pla_top/N59 ;
   wire \pla_top/instruction_valid ;
   wire \addr_calc/N224 ;
   wire \addr_calc/N223 ;
   wire \addr_calc/N220 ;
   wire \addr_calc/N219 ;
   wire \addr_calc/N217 ;
   wire \addr_calc/N216 ;
   wire \addr_calc/iir_write_addr[31] ;
   wire \addr_calc/iir_write_addr[30] ;
   wire \addr_calc/iir_write_addr[29] ;
   wire \addr_calc/iir_write_addr[28] ;
   wire \addr_calc/iir_write_addr[27] ;
   wire \addr_calc/iir_write_addr[26] ;
   wire \addr_calc/iir_write_addr[24] ;
   wire \addr_calc/iir_write_addr[23] ;
   wire \addr_calc/iir_write_addr[22] ;
   wire \addr_calc/iir_write_addr[20] ;
   wire \addr_calc/iir_write_addr[18] ;
   wire \addr_calc/iir_write_addr[17] ;
   wire \addr_calc/iir_write_addr[15] ;
   wire \addr_calc/iir_write_addr[14] ;
   wire \addr_calc/iir_write_addr[13] ;
   wire \addr_calc/iir_write_addr[12] ;
   wire \addr_calc/iir_write_addr[11] ;
   wire \addr_calc/iir_write_addr[8] ;
   wire \addr_calc/iir_write_addr[7] ;
   wire \addr_calc/iir_write_addr[6] ;
   wire \addr_calc/iir_write_addr[5] ;
   wire \addr_calc/iir_write_addr[4] ;
   wire \addr_calc/iir_write_addr[3] ;
   wire \addr_calc/iir_write_addr[2] ;
   wire \addr_calc/iir_write_addr[1] ;
   wire \addr_calc/iir_write_addr[0] ;
   wire \addr_calc/iir_read_addr[31] ;
   wire \addr_calc/iir_read_addr[30] ;
   wire \addr_calc/iir_read_addr[29] ;
   wire \addr_calc/iir_read_addr[28] ;
   wire \addr_calc/iir_read_addr[27] ;
   wire \addr_calc/iir_read_addr[26] ;
   wire \addr_calc/iir_read_addr[25] ;
   wire \addr_calc/iir_read_addr[23] ;
   wire \addr_calc/iir_read_addr[22] ;
   wire \addr_calc/iir_read_addr[21] ;
   wire \addr_calc/iir_read_addr[20] ;
   wire \addr_calc/iir_read_addr[19] ;
   wire \addr_calc/iir_read_addr[18] ;
   wire \addr_calc/iir_read_addr[17] ;
   wire \addr_calc/iir_read_addr[16] ;
   wire \addr_calc/iir_read_addr[14] ;
   wire \addr_calc/iir_read_addr[13] ;
   wire \addr_calc/iir_read_addr[12] ;
   wire \addr_calc/iir_read_addr[11] ;
   wire \addr_calc/iir_read_addr[10] ;
   wire \addr_calc/iir_read_addr[8] ;
   wire \addr_calc/iir_read_addr[7] ;
   wire \addr_calc/iir_read_addr[6] ;
   wire \addr_calc/iir_read_addr[5] ;
   wire \addr_calc/iir_read_addr[4] ;
   wire \addr_calc/iir_read_addr[3] ;
   wire \addr_calc/iir_read_addr[2] ;
   wire \addr_calc/iir_read_addr[1] ;
   wire \addr_calc/iir_read_addr[0] ;
   wire \addr_calc/fir_write_addr[31] ;
   wire \addr_calc/fir_write_addr[30] ;
   wire \addr_calc/fir_write_addr[29] ;
   wire \addr_calc/fir_write_addr[28] ;
   wire \addr_calc/fir_write_addr[27] ;
   wire \addr_calc/fir_write_addr[26] ;
   wire \addr_calc/fir_write_addr[25] ;
   wire \addr_calc/fir_write_addr[24] ;
   wire \addr_calc/fir_write_addr[23] ;
   wire \addr_calc/fir_write_addr[22] ;
   wire \addr_calc/fir_write_addr[21] ;
   wire \addr_calc/fir_write_addr[20] ;
   wire \addr_calc/fir_write_addr[19] ;
   wire \addr_calc/fir_write_addr[18] ;
   wire \addr_calc/fir_write_addr[17] ;
   wire \addr_calc/fir_write_addr[16] ;
   wire \addr_calc/fir_write_addr[15] ;
   wire \addr_calc/fir_write_addr[14] ;
   wire \addr_calc/fir_write_addr[13] ;
   wire \addr_calc/fir_write_addr[12] ;
   wire \addr_calc/fir_write_addr[11] ;
   wire \addr_calc/fir_write_addr[10] ;
   wire \addr_calc/fir_write_addr[9] ;
   wire \addr_calc/fir_write_addr[8] ;
   wire \addr_calc/fir_write_addr[7] ;
   wire \addr_calc/fir_write_addr[6] ;
   wire \addr_calc/fir_write_addr[5] ;
   wire \addr_calc/fir_write_addr[4] ;
   wire \addr_calc/fir_write_addr[3] ;
   wire \addr_calc/fir_write_addr[2] ;
   wire \addr_calc/fir_write_addr[1] ;
   wire \addr_calc/fir_write_addr[0] ;
   wire \addr_calc/fir_read_addr[31] ;
   wire \addr_calc/fir_read_addr[30] ;
   wire \addr_calc/fir_read_addr[29] ;
   wire \addr_calc/fir_read_addr[28] ;
   wire \addr_calc/fir_read_addr[27] ;
   wire \addr_calc/fir_read_addr[26] ;
   wire \addr_calc/fir_read_addr[25] ;
   wire \addr_calc/fir_read_addr[24] ;
   wire \addr_calc/fir_read_addr[23] ;
   wire \addr_calc/fir_read_addr[22] ;
   wire \addr_calc/fir_read_addr[21] ;
   wire \addr_calc/fir_read_addr[20] ;
   wire \addr_calc/fir_read_addr[19] ;
   wire \addr_calc/fir_read_addr[18] ;
   wire \addr_calc/fir_read_addr[17] ;
   wire \addr_calc/fir_read_addr[16] ;
   wire \addr_calc/fir_read_addr[15] ;
   wire \addr_calc/fir_read_addr[14] ;
   wire \addr_calc/fir_read_addr[13] ;
   wire \addr_calc/fir_read_addr[12] ;
   wire \addr_calc/fir_read_addr[11] ;
   wire \addr_calc/fir_read_addr[10] ;
   wire \addr_calc/fir_read_addr[9] ;
   wire \addr_calc/fir_read_addr[8] ;
   wire \addr_calc/fir_read_addr[7] ;
   wire \addr_calc/fir_read_addr[6] ;
   wire \addr_calc/fir_read_addr[5] ;
   wire \addr_calc/fir_read_addr[4] ;
   wire \addr_calc/fir_read_addr[3] ;
   wire \addr_calc/fir_read_addr[2] ;
   wire \addr_calc/fir_read_addr[1] ;
   wire \addr_calc/fir_read_addr[0] ;
   wire \addr_calc/fft_write_addr[31] ;
   wire \addr_calc/fft_write_addr[30] ;
   wire \addr_calc/fft_write_addr[29] ;
   wire \addr_calc/fft_write_addr[28] ;
   wire \addr_calc/fft_write_addr[27] ;
   wire \addr_calc/fft_write_addr[26] ;
   wire \addr_calc/fft_write_addr[25] ;
   wire \addr_calc/fft_write_addr[24] ;
   wire \addr_calc/fft_write_addr[23] ;
   wire \addr_calc/fft_write_addr[22] ;
   wire \addr_calc/fft_write_addr[21] ;
   wire \addr_calc/fft_write_addr[20] ;
   wire \addr_calc/fft_write_addr[19] ;
   wire \addr_calc/fft_write_addr[18] ;
   wire \addr_calc/fft_write_addr[17] ;
   wire \addr_calc/fft_write_addr[16] ;
   wire \addr_calc/fft_write_addr[15] ;
   wire \addr_calc/fft_write_addr[14] ;
   wire \addr_calc/fft_write_addr[13] ;
   wire \addr_calc/fft_write_addr[12] ;
   wire \addr_calc/fft_write_addr[11] ;
   wire \addr_calc/fft_write_addr[10] ;
   wire \addr_calc/fft_write_addr[9] ;
   wire \addr_calc/fft_write_addr[8] ;
   wire \addr_calc/fft_write_addr[7] ;
   wire \addr_calc/fft_write_addr[6] ;
   wire \addr_calc/fft_write_addr[5] ;
   wire \addr_calc/fft_write_addr[4] ;
   wire \addr_calc/fft_write_addr[3] ;
   wire \addr_calc/fft_write_addr[2] ;
   wire \addr_calc/fft_write_addr[1] ;
   wire \addr_calc/fft_write_addr[0] ;
   wire \addr_calc/fft_read_addr[31] ;
   wire \addr_calc/fft_read_addr[27] ;
   wire \addr_calc/fft_read_addr[26] ;
   wire \addr_calc/fft_read_addr[25] ;
   wire \addr_calc/fft_read_addr[24] ;
   wire \addr_calc/fft_read_addr[23] ;
   wire \addr_calc/fft_read_addr[22] ;
   wire \addr_calc/fft_read_addr[21] ;
   wire \addr_calc/fft_read_addr[20] ;
   wire \addr_calc/fft_read_addr[19] ;
   wire \addr_calc/fft_read_addr[18] ;
   wire \addr_calc/fft_read_addr[17] ;
   wire \addr_calc/fft_read_addr[16] ;
   wire \addr_calc/fft_read_addr[15] ;
   wire \addr_calc/fft_read_addr[14] ;
   wire \addr_calc/fft_read_addr[13] ;
   wire \addr_calc/fft_read_addr[12] ;
   wire \addr_calc/fft_read_addr[11] ;
   wire \addr_calc/fft_read_addr[10] ;
   wire \addr_calc/fft_read_addr[9] ;
   wire \addr_calc/fft_read_addr[8] ;
   wire \addr_calc/fft_read_addr[7] ;
   wire \addr_calc/fft_read_addr[6] ;
   wire \addr_calc/fft_read_addr[5] ;
   wire \addr_calc/fft_read_addr[4] ;
   wire \addr_calc/fft_read_addr[3] ;
   wire \addr_calc/fft_read_addr[2] ;
   wire \addr_calc/fft_read_addr[1] ;
   wire \addr_calc/fft_read_addr[0] ;
   wire \addr_calc/N191 ;
   wire \addr_calc/N159 ;
   wire \addr_calc/N99 ;
   wire \addr_calc/N95 ;
   wire \addr_calc/N63 ;
   wire \addr_calc/N9 ;
   wire \data_cntl/N267 ;
   wire \data_cntl/N266 ;
   wire \data_cntl/N265 ;
   wire \data_cntl/N264 ;
   wire \data_cntl/N263 ;
   wire \data_cntl/N262 ;
   wire \data_cntl/N261 ;
   wire \data_cntl/N260 ;
   wire \data_cntl/N259 ;
   wire \data_cntl/N258 ;
   wire \data_cntl/N257 ;
   wire \data_cntl/N256 ;
   wire \data_cntl/N255 ;
   wire \data_cntl/N254 ;
   wire \data_cntl/N253 ;
   wire \data_cntl/N252 ;
   wire \data_cntl/N251 ;
   wire \data_cntl/N250 ;
   wire \data_cntl/N191 ;
   wire \data_cntl/N159 ;
   wire \data_cntl/N99 ;
   wire \data_cntl/N95 ;
   wire \data_cntl/N63 ;
   wire \data_cntl/N9 ;
   wire \addr_calc/fft_read_calc/count[31] ;
   wire \addr_calc/fft_read_calc/count[30] ;
   wire \addr_calc/fft_read_calc/count[29] ;
   wire \addr_calc/fft_read_calc/count[28] ;
   wire \addr_calc/fft_read_calc/count[27] ;
   wire \addr_calc/fft_read_calc/count[26] ;
   wire \addr_calc/fft_read_calc/count[25] ;
   wire \addr_calc/fft_read_calc/count[24] ;
   wire \addr_calc/fft_read_calc/count[23] ;
   wire \addr_calc/fft_read_calc/count[22] ;
   wire \addr_calc/fft_read_calc/count[21] ;
   wire \addr_calc/fft_read_calc/count[20] ;
   wire \addr_calc/fft_read_calc/count[19] ;
   wire \addr_calc/fft_read_calc/count[18] ;
   wire \addr_calc/fft_read_calc/count[17] ;
   wire \addr_calc/fft_read_calc/count[16] ;
   wire \addr_calc/fft_read_calc/count[15] ;
   wire \addr_calc/fft_read_calc/count[14] ;
   wire \addr_calc/fft_read_calc/count[13] ;
   wire \addr_calc/fft_read_calc/count[12] ;
   wire \addr_calc/fft_read_calc/count[11] ;
   wire \addr_calc/fft_read_calc/count[10] ;
   wire \addr_calc/fft_read_calc/count[9] ;
   wire \addr_calc/fft_read_calc/count[8] ;
   wire \addr_calc/fft_read_calc/count[7] ;
   wire \addr_calc/fft_read_calc/count[6] ;
   wire \addr_calc/fft_read_calc/count[5] ;
   wire \addr_calc/fft_read_calc/count[4] ;
   wire \addr_calc/fft_read_calc/count[3] ;
   wire \addr_calc/fft_read_calc/count[2] ;
   wire \addr_calc/fft_read_calc/count[1] ;
   wire \addr_calc/fft_read_calc/count[0] ;
   wire \addr_calc/fft_write_calc/count[31] ;
   wire \addr_calc/fft_write_calc/count[30] ;
   wire \addr_calc/fft_write_calc/count[29] ;
   wire \addr_calc/fft_write_calc/count[28] ;
   wire \addr_calc/fft_write_calc/count[27] ;
   wire \addr_calc/fft_write_calc/count[26] ;
   wire \addr_calc/fft_write_calc/count[25] ;
   wire \addr_calc/fft_write_calc/count[24] ;
   wire \addr_calc/fft_write_calc/count[23] ;
   wire \addr_calc/fft_write_calc/count[22] ;
   wire \addr_calc/fft_write_calc/count[21] ;
   wire \addr_calc/fft_write_calc/count[20] ;
   wire \addr_calc/fft_write_calc/count[19] ;
   wire \addr_calc/fft_write_calc/count[18] ;
   wire \addr_calc/fft_write_calc/count[17] ;
   wire \addr_calc/fft_write_calc/count[16] ;
   wire \addr_calc/fft_write_calc/count[15] ;
   wire \addr_calc/fft_write_calc/count[14] ;
   wire \addr_calc/fft_write_calc/count[13] ;
   wire \addr_calc/fft_write_calc/count[12] ;
   wire \addr_calc/fft_write_calc/count[11] ;
   wire \addr_calc/fft_write_calc/count[10] ;
   wire \addr_calc/fft_write_calc/count[9] ;
   wire \addr_calc/fft_write_calc/count[8] ;
   wire \addr_calc/fft_write_calc/count[7] ;
   wire \addr_calc/fft_write_calc/count[6] ;
   wire \addr_calc/fft_write_calc/count[5] ;
   wire \addr_calc/fft_write_calc/count[4] ;
   wire \addr_calc/fft_write_calc/count[3] ;
   wire \addr_calc/fft_write_calc/count[2] ;
   wire \addr_calc/fft_write_calc/count[1] ;
   wire \addr_calc/fft_write_calc/count[0] ;
   wire \addr_calc/fir_read_calc/count[31] ;
   wire \addr_calc/fir_read_calc/count[30] ;
   wire \addr_calc/fir_read_calc/count[29] ;
   wire \addr_calc/fir_read_calc/count[28] ;
   wire \addr_calc/fir_read_calc/count[27] ;
   wire \addr_calc/fir_read_calc/count[26] ;
   wire \addr_calc/fir_read_calc/count[25] ;
   wire \addr_calc/fir_read_calc/count[24] ;
   wire \addr_calc/fir_read_calc/count[23] ;
   wire \addr_calc/fir_read_calc/count[22] ;
   wire \addr_calc/fir_read_calc/count[21] ;
   wire \addr_calc/fir_read_calc/count[20] ;
   wire \addr_calc/fir_read_calc/count[19] ;
   wire \addr_calc/fir_read_calc/count[18] ;
   wire \addr_calc/fir_read_calc/count[17] ;
   wire \addr_calc/fir_read_calc/count[16] ;
   wire \addr_calc/fir_read_calc/count[15] ;
   wire \addr_calc/fir_read_calc/count[14] ;
   wire \addr_calc/fir_read_calc/count[13] ;
   wire \addr_calc/fir_read_calc/count[12] ;
   wire \addr_calc/fir_read_calc/count[11] ;
   wire \addr_calc/fir_read_calc/count[10] ;
   wire \addr_calc/fir_read_calc/count[9] ;
   wire \addr_calc/fir_read_calc/count[8] ;
   wire \addr_calc/fir_read_calc/count[7] ;
   wire \addr_calc/fir_read_calc/count[6] ;
   wire \addr_calc/fir_read_calc/count[5] ;
   wire \addr_calc/fir_read_calc/count[4] ;
   wire \addr_calc/fir_read_calc/count[3] ;
   wire \addr_calc/fir_read_calc/count[2] ;
   wire \addr_calc/fir_read_calc/count[1] ;
   wire \addr_calc/fir_read_calc/count[0] ;
   wire \addr_calc/fir_write_calc/count[31] ;
   wire \addr_calc/fir_write_calc/count[30] ;
   wire \addr_calc/fir_write_calc/count[29] ;
   wire \addr_calc/fir_write_calc/count[28] ;
   wire \addr_calc/fir_write_calc/count[27] ;
   wire \addr_calc/fir_write_calc/count[26] ;
   wire \addr_calc/fir_write_calc/count[25] ;
   wire \addr_calc/fir_write_calc/count[24] ;
   wire \addr_calc/fir_write_calc/count[23] ;
   wire \addr_calc/fir_write_calc/count[22] ;
   wire \addr_calc/fir_write_calc/count[21] ;
   wire \addr_calc/fir_write_calc/count[20] ;
   wire \addr_calc/fir_write_calc/count[19] ;
   wire \addr_calc/fir_write_calc/count[18] ;
   wire \addr_calc/fir_write_calc/count[17] ;
   wire \addr_calc/fir_write_calc/count[16] ;
   wire \addr_calc/fir_write_calc/count[15] ;
   wire \addr_calc/fir_write_calc/count[14] ;
   wire \addr_calc/fir_write_calc/count[13] ;
   wire \addr_calc/fir_write_calc/count[12] ;
   wire \addr_calc/fir_write_calc/count[11] ;
   wire \addr_calc/fir_write_calc/count[10] ;
   wire \addr_calc/fir_write_calc/count[9] ;
   wire \addr_calc/fir_write_calc/count[8] ;
   wire \addr_calc/fir_write_calc/count[7] ;
   wire \addr_calc/fir_write_calc/count[6] ;
   wire \addr_calc/fir_write_calc/count[5] ;
   wire \addr_calc/fir_write_calc/count[4] ;
   wire \addr_calc/fir_write_calc/count[3] ;
   wire \addr_calc/fir_write_calc/count[2] ;
   wire \addr_calc/fir_write_calc/count[1] ;
   wire \addr_calc/fir_write_calc/count[0] ;
   wire \addr_calc/iir_read_calc/count[31] ;
   wire \addr_calc/iir_read_calc/count[30] ;
   wire \addr_calc/iir_read_calc/count[29] ;
   wire \addr_calc/iir_read_calc/count[28] ;
   wire \addr_calc/iir_read_calc/count[27] ;
   wire \addr_calc/iir_read_calc/count[26] ;
   wire \addr_calc/iir_read_calc/count[25] ;
   wire \addr_calc/iir_read_calc/count[24] ;
   wire \addr_calc/iir_read_calc/count[23] ;
   wire \addr_calc/iir_read_calc/count[22] ;
   wire \addr_calc/iir_read_calc/count[21] ;
   wire \addr_calc/iir_read_calc/count[20] ;
   wire \addr_calc/iir_read_calc/count[19] ;
   wire \addr_calc/iir_read_calc/count[18] ;
   wire \addr_calc/iir_read_calc/count[17] ;
   wire \addr_calc/iir_read_calc/count[16] ;
   wire \addr_calc/iir_read_calc/count[15] ;
   wire \addr_calc/iir_read_calc/count[14] ;
   wire \addr_calc/iir_read_calc/count[13] ;
   wire \addr_calc/iir_read_calc/count[12] ;
   wire \addr_calc/iir_read_calc/count[11] ;
   wire \addr_calc/iir_read_calc/count[10] ;
   wire \addr_calc/iir_read_calc/count[9] ;
   wire \addr_calc/iir_read_calc/count[8] ;
   wire \addr_calc/iir_read_calc/count[7] ;
   wire \addr_calc/iir_read_calc/count[6] ;
   wire \addr_calc/iir_read_calc/count[5] ;
   wire \addr_calc/iir_read_calc/count[4] ;
   wire \addr_calc/iir_read_calc/count[3] ;
   wire \addr_calc/iir_read_calc/count[2] ;
   wire \addr_calc/iir_read_calc/count[1] ;
   wire \addr_calc/iir_read_calc/count[0] ;
   wire \addr_calc/iir_write_calc/count[31] ;
   wire \addr_calc/iir_write_calc/count[30] ;
   wire \addr_calc/iir_write_calc/count[29] ;
   wire \addr_calc/iir_write_calc/count[28] ;
   wire \addr_calc/iir_write_calc/count[27] ;
   wire \addr_calc/iir_write_calc/count[26] ;
   wire \addr_calc/iir_write_calc/count[25] ;
   wire \addr_calc/iir_write_calc/count[24] ;
   wire \addr_calc/iir_write_calc/count[23] ;
   wire \addr_calc/iir_write_calc/count[22] ;
   wire \addr_calc/iir_write_calc/count[21] ;
   wire \addr_calc/iir_write_calc/count[20] ;
   wire \addr_calc/iir_write_calc/count[19] ;
   wire \addr_calc/iir_write_calc/count[18] ;
   wire \addr_calc/iir_write_calc/count[17] ;
   wire \addr_calc/iir_write_calc/count[16] ;
   wire \addr_calc/iir_write_calc/count[15] ;
   wire \addr_calc/iir_write_calc/count[14] ;
   wire \addr_calc/iir_write_calc/count[13] ;
   wire \addr_calc/iir_write_calc/count[12] ;
   wire \addr_calc/iir_write_calc/count[11] ;
   wire \addr_calc/iir_write_calc/count[10] ;
   wire \addr_calc/iir_write_calc/count[9] ;
   wire \addr_calc/iir_write_calc/count[8] ;
   wire \addr_calc/iir_write_calc/count[7] ;
   wire \addr_calc/iir_write_calc/count[6] ;
   wire \addr_calc/iir_write_calc/count[5] ;
   wire \addr_calc/iir_write_calc/count[4] ;
   wire \addr_calc/iir_write_calc/count[3] ;
   wire \addr_calc/iir_write_calc/count[2] ;
   wire \addr_calc/iir_write_calc/count[1] ;
   wire \addr_calc/iir_write_calc/count[0] ;
   wire \addr_calc/fft_read_calc/counter/N73 ;
   wire \addr_calc/fft_read_calc/counter/N72 ;
   wire \addr_calc/fft_read_calc/counter/N71 ;
   wire \addr_calc/fft_read_calc/counter/N70 ;
   wire \addr_calc/fft_read_calc/counter/N68 ;
   wire \addr_calc/fft_read_calc/counter/N67 ;
   wire \addr_calc/fft_read_calc/counter/N66 ;
   wire \addr_calc/fft_read_calc/counter/N65 ;
   wire \addr_calc/fft_read_calc/counter/N63 ;
   wire \addr_calc/fft_read_calc/counter/N62 ;
   wire \addr_calc/fft_read_calc/counter/N58 ;
   wire \addr_calc/fft_read_calc/counter/N57 ;
   wire \addr_calc/fft_read_calc/counter/N56 ;
   wire \addr_calc/fft_read_calc/counter/N55 ;
   wire \addr_calc/fft_read_calc/counter/N53 ;
   wire \addr_calc/fft_read_calc/counter/N52 ;
   wire \addr_calc/fft_read_calc/counter/N51 ;
   wire \addr_calc/fft_read_calc/counter/N50 ;
   wire \addr_calc/fft_read_calc/counter/N48 ;
   wire \addr_calc/fft_read_calc/counter/N46 ;
   wire \addr_calc/fft_read_calc/counter/N45 ;
   wire \addr_calc/fft_read_calc/counter/N44 ;
   wire \addr_calc/fft_read_calc/counter/N38 ;
   wire \addr_calc/fft_write_calc/counter/N74 ;
   wire \addr_calc/fft_write_calc/counter/N73 ;
   wire \addr_calc/fft_write_calc/counter/N72 ;
   wire \addr_calc/fft_write_calc/counter/N71 ;
   wire \addr_calc/fft_write_calc/counter/N68 ;
   wire \addr_calc/fft_write_calc/counter/N66 ;
   wire \addr_calc/fft_write_calc/counter/N64 ;
   wire \addr_calc/fft_write_calc/counter/N62 ;
   wire \addr_calc/fft_write_calc/counter/N60 ;
   wire \addr_calc/fft_write_calc/counter/N59 ;
   wire \addr_calc/fft_write_calc/counter/N58 ;
   wire \addr_calc/fft_write_calc/counter/N57 ;
   wire \addr_calc/fft_write_calc/counter/N56 ;
   wire \addr_calc/fft_write_calc/counter/N55 ;
   wire \addr_calc/fft_write_calc/counter/N53 ;
   wire \addr_calc/fft_write_calc/counter/N52 ;
   wire \addr_calc/fft_write_calc/counter/N51 ;
   wire \addr_calc/fft_write_calc/counter/N50 ;
   wire \addr_calc/fft_write_calc/counter/N47 ;
   wire \addr_calc/fft_write_calc/counter/N46 ;
   wire \addr_calc/fft_write_calc/counter/N43 ;
   wire \addr_calc/fft_write_calc/counter/N38 ;
   wire \addr_calc/fir_read_calc/counter/N73 ;
   wire \addr_calc/fir_read_calc/counter/N72 ;
   wire \addr_calc/fir_read_calc/counter/N71 ;
   wire \addr_calc/fir_read_calc/counter/N67 ;
   wire \addr_calc/fir_read_calc/counter/N66 ;
   wire \addr_calc/fir_read_calc/counter/N65 ;
   wire \addr_calc/fir_read_calc/counter/N64 ;
   wire \addr_calc/fir_read_calc/counter/N63 ;
   wire \addr_calc/fir_read_calc/counter/N62 ;
   wire \addr_calc/fir_read_calc/counter/N61 ;
   wire \addr_calc/fir_read_calc/counter/N60 ;
   wire \addr_calc/fir_read_calc/counter/N59 ;
   wire \addr_calc/fir_read_calc/counter/N57 ;
   wire \addr_calc/fir_read_calc/counter/N56 ;
   wire \addr_calc/fir_read_calc/counter/N55 ;
   wire \addr_calc/fir_read_calc/counter/N54 ;
   wire \addr_calc/fir_read_calc/counter/N53 ;
   wire \addr_calc/fir_read_calc/counter/N52 ;
   wire \addr_calc/fir_read_calc/counter/N51 ;
   wire \addr_calc/fir_read_calc/counter/N50 ;
   wire \addr_calc/fir_read_calc/counter/N49 ;
   wire \addr_calc/fir_read_calc/counter/N48 ;
   wire \addr_calc/fir_read_calc/counter/N47 ;
   wire \addr_calc/fir_read_calc/counter/N45 ;
   wire \addr_calc/fir_read_calc/counter/N44 ;
   wire \addr_calc/fir_read_calc/counter/N38 ;
   wire \addr_calc/fir_write_calc/counter/N74 ;
   wire \addr_calc/fir_write_calc/counter/N73 ;
   wire \addr_calc/fir_write_calc/counter/N72 ;
   wire \addr_calc/fir_write_calc/counter/N71 ;
   wire \addr_calc/fir_write_calc/counter/N70 ;
   wire \addr_calc/fir_write_calc/counter/N68 ;
   wire \addr_calc/fir_write_calc/counter/N67 ;
   wire \addr_calc/fir_write_calc/counter/N66 ;
   wire \addr_calc/fir_write_calc/counter/N65 ;
   wire \addr_calc/fir_write_calc/counter/N62 ;
   wire \addr_calc/fir_write_calc/counter/N61 ;
   wire \addr_calc/fir_write_calc/counter/N60 ;
   wire \addr_calc/fir_write_calc/counter/N59 ;
   wire \addr_calc/fir_write_calc/counter/N57 ;
   wire \addr_calc/fir_write_calc/counter/N56 ;
   wire \addr_calc/fir_write_calc/counter/N54 ;
   wire \addr_calc/fir_write_calc/counter/N52 ;
   wire \addr_calc/fir_write_calc/counter/N51 ;
   wire \addr_calc/fir_write_calc/counter/N49 ;
   wire \addr_calc/fir_write_calc/counter/N48 ;
   wire \addr_calc/fir_write_calc/counter/N46 ;
   wire \addr_calc/fir_write_calc/counter/N45 ;
   wire \addr_calc/fir_write_calc/counter/N43 ;
   wire \addr_calc/fir_write_calc/counter/N38 ;
   wire \addr_calc/iir_read_calc/counter/N74 ;
   wire \addr_calc/iir_read_calc/counter/N73 ;
   wire \addr_calc/iir_read_calc/counter/N72 ;
   wire \addr_calc/iir_read_calc/counter/N71 ;
   wire \addr_calc/iir_read_calc/counter/N68 ;
   wire \addr_calc/iir_read_calc/counter/N67 ;
   wire \addr_calc/iir_read_calc/counter/N63 ;
   wire \addr_calc/iir_read_calc/counter/N62 ;
   wire \addr_calc/iir_read_calc/counter/N61 ;
   wire \addr_calc/iir_read_calc/counter/N60 ;
   wire \addr_calc/iir_read_calc/counter/N59 ;
   wire \addr_calc/iir_read_calc/counter/N58 ;
   wire \addr_calc/iir_read_calc/counter/N57 ;
   wire \addr_calc/iir_read_calc/counter/N55 ;
   wire \addr_calc/iir_read_calc/counter/N54 ;
   wire \addr_calc/iir_read_calc/counter/N53 ;
   wire \addr_calc/iir_read_calc/counter/N52 ;
   wire \addr_calc/iir_read_calc/counter/N51 ;
   wire \addr_calc/iir_read_calc/counter/N50 ;
   wire \addr_calc/iir_read_calc/counter/N48 ;
   wire \addr_calc/iir_read_calc/counter/N46 ;
   wire \addr_calc/iir_read_calc/counter/N45 ;
   wire \addr_calc/iir_read_calc/counter/N44 ;
   wire \addr_calc/iir_write_calc/counter/N74 ;
   wire \addr_calc/iir_write_calc/counter/N73 ;
   wire \addr_calc/iir_write_calc/counter/N72 ;
   wire \addr_calc/iir_write_calc/counter/N71 ;
   wire \addr_calc/iir_write_calc/counter/N70 ;
   wire \addr_calc/iir_write_calc/counter/N69 ;
   wire \addr_calc/iir_write_calc/counter/N68 ;
   wire \addr_calc/iir_write_calc/counter/N67 ;
   wire \addr_calc/iir_write_calc/counter/N66 ;
   wire \addr_calc/iir_write_calc/counter/N65 ;
   wire \addr_calc/iir_write_calc/counter/N62 ;
   wire \addr_calc/iir_write_calc/counter/N60 ;
   wire \addr_calc/iir_write_calc/counter/N57 ;
   wire \addr_calc/iir_write_calc/counter/N56 ;
   wire \addr_calc/iir_write_calc/counter/N55 ;
   wire \addr_calc/iir_write_calc/counter/N54 ;
   wire \addr_calc/iir_write_calc/counter/N53 ;
   wire \addr_calc/iir_write_calc/counter/N52 ;
   wire \addr_calc/iir_write_calc/counter/N51 ;
   wire \addr_calc/iir_write_calc/counter/N50 ;
   wire \addr_calc/iir_write_calc/counter/N49 ;
   wire \addr_calc/iir_write_calc/counter/N48 ;
   wire \addr_calc/iir_write_calc/counter/N47 ;
   wire \addr_calc/iir_write_calc/counter/N46 ;
   wire \addr_calc/iir_write_calc/counter/N45 ;
   wire \addr_calc/iir_write_calc/counter/N44 ;
   wire n3;
   wire n67;
   wire n131;
   wire n195;
   wire n259;
   wire n323;
   wire n387;
   wire n451;
   wire n515;
   wire n579;
   wire n643;
   wire n707;
   wire n783;
   wire n785;
   wire n787;
   wire n790;
   wire n791;
   wire n792;
   wire n793;
   wire n795;
   wire n796;
   wire n797;
   wire n798;
   wire n801;
   wire n802;
   wire n810;
   wire n811;
   wire n812;
   wire n813;
   wire n814;
   wire n815;
   wire n816;
   wire n817;
   wire n828;
   wire n829;
   wire n830;
   wire n831;
   wire n832;
   wire n833;
   wire n842;
   wire n843;
   wire n844;
   wire n845;
   wire n846;
   wire n847;
   wire n861;
   wire n862;
   wire n863;
   wire n864;
   wire n865;
   wire n866;
   wire n867;
   wire n868;
   wire n869;
   wire n870;
   wire n871;
   wire n872;
   wire n873;
   wire n876;
   wire n877;
   wire n878;
   wire n879;
   wire n880;
   wire n881;
   wire n882;
   wire n883;
   wire n884;
   wire n885;
   wire n886;
   wire n887;
   wire n888;
   wire n889;
   wire n890;
   wire n891;
   wire n892;
   wire n893;
   wire n894;
   wire n895;
   wire n897;
   wire n898;
   wire n899;
   wire n900;
   wire n901;
   wire n902;
   wire n903;
   wire n904;
   wire n905;
   wire n906;
   wire n907;
   wire n908;
   wire n915;
   wire n916;
   wire n917;
   wire n918;
   wire n919;
   wire n920;
   wire n921;
   wire n922;
   wire n923;
   wire n924;
   wire n925;
   wire n926;
   wire n927;
   wire n928;
   wire n929;
   wire n930;
   wire n931;
   wire n932;
   wire n933;
   wire n934;
   wire n935;
   wire n936;
   wire n937;
   wire n938;
   wire n939;
   wire n940;
   wire n941;
   wire n942;
   wire n943;
   wire n944;
   wire n945;
   wire n946;
   wire n947;
   wire n948;
   wire n949;
   wire n950;
   wire n951;
   wire n952;
   wire n953;
   wire n954;
   wire n955;
   wire n956;
   wire n957;
   wire n958;
   wire n959;
   wire n960;
   wire n961;
   wire n962;
   wire n963;
   wire n964;
   wire n965;
   wire n966;
   wire n967;
   wire n968;
   wire n969;
   wire n970;
   wire n971;
   wire n972;
   wire n973;
   wire n974;
   wire n975;
   wire n976;
   wire n977;
   wire n978;
   wire n979;
   wire n980;
   wire n981;
   wire n982;
   wire n983;
   wire n984;
   wire n985;
   wire n986;
   wire n987;
   wire n988;
   wire n989;
   wire n990;
   wire n991;
   wire n992;
   wire n993;
   wire n994;
   wire n995;
   wire n996;
   wire n997;
   wire n998;
   wire n999;
   wire n1000;
   wire n1001;
   wire n1002;
   wire n1003;
   wire n1004;
   wire n1005;
   wire n1006;
   wire n1007;
   wire n1008;
   wire n1009;
   wire n1010;
   wire n1011;
   wire n1012;
   wire n1013;
   wire n1014;
   wire n1015;
   wire n1016;
   wire n1017;
   wire n1018;
   wire n1019;
   wire n1020;
   wire n1021;
   wire n1022;
   wire n1023;
   wire n1024;
   wire n1025;
   wire n1026;
   wire n1027;
   wire n1028;
   wire n1029;
   wire n1030;
   wire n1031;
   wire n1032;
   wire n1033;
   wire n1034;
   wire n1035;
   wire n1036;
   wire n1037;
   wire n1038;
   wire n1039;
   wire n1040;
   wire n1041;
   wire n1042;
   wire n1043;
   wire n1044;
   wire n1045;
   wire n1046;
   wire n1047;
   wire n1048;
   wire n1049;
   wire n1050;
   wire n1051;
   wire n1052;
   wire n1053;
   wire n1054;
   wire n1055;
   wire n1056;
   wire n1057;
   wire n1058;
   wire n1059;
   wire n1060;
   wire n1061;
   wire n1062;
   wire n1063;
   wire n1064;
   wire n1065;
   wire n1066;
   wire n1067;
   wire n1068;
   wire n1069;
   wire n1070;
   wire n1071;
   wire n1072;
   wire n1073;
   wire n1074;
   wire n1075;
   wire n1076;
   wire n1077;
   wire n1078;
   wire n1079;
   wire n1080;
   wire n1081;
   wire n1082;
   wire n1083;
   wire n1084;
   wire n1085;
   wire n1086;
   wire n1087;
   wire n1088;
   wire n1089;
   wire n1090;
   wire n1091;
   wire n1092;
   wire n1093;
   wire n1094;
   wire n1095;
   wire n1096;
   wire n1097;
   wire n1098;
   wire n1099;
   wire n1100;
   wire n1101;
   wire n1102;
   wire n1103;
   wire n1104;
   wire n1105;
   wire n1106;
   wire n1107;
   wire n1108;
   wire n1109;
   wire n1110;
   wire n1111;
   wire n1112;
   wire n1113;
   wire n1114;
   wire n1115;
   wire n1116;
   wire n1117;
   wire n1118;
   wire n1119;
   wire n1120;
   wire n1121;
   wire n1122;
   wire n1123;
   wire n1124;
   wire n1125;
   wire n1126;
   wire n1127;
   wire n1128;
   wire n1129;
   wire n1130;
   wire n1131;
   wire n1132;
   wire n1133;
   wire n1134;
   wire n1135;
   wire n1136;
   wire \add_x_19_4/n222 ;
   wire \add_x_19_4/n221 ;
   wire \add_x_19_4/n219 ;
   wire \add_x_19_4/n217 ;
   wire \add_x_19_4/n213 ;
   wire \add_x_19_4/n212 ;
   wire \add_x_19_4/n207 ;
   wire \add_x_19_4/n206 ;
   wire \add_x_19_4/n204 ;
   wire \add_x_19_4/n202 ;
   wire \add_x_19_4/n199 ;
   wire \add_x_19_4/n196 ;
   wire \add_x_19_4/n191 ;
   wire \add_x_19_4/n189 ;
   wire \add_x_19_4/n188 ;
   wire \add_x_19_4/n187 ;
   wire \add_x_19_4/n186 ;
   wire \add_x_19_4/n185 ;
   wire \add_x_19_4/n184 ;
   wire \add_x_19_4/n182 ;
   wire \add_x_19_4/n181 ;
   wire \add_x_19_4/n178 ;
   wire \add_x_19_4/n176 ;
   wire \add_x_19_4/n175 ;
   wire \add_x_19_4/n171 ;
   wire \add_x_19_4/n170 ;
   wire \add_x_19_4/n169 ;
   wire \add_x_19_4/n168 ;
   wire \add_x_19_4/n167 ;
   wire \add_x_19_4/n166 ;
   wire \add_x_19_4/n165 ;
   wire \add_x_19_4/n163 ;
   wire \add_x_19_4/n162 ;
   wire \add_x_19_4/n160 ;
   wire \add_x_19_4/n157 ;
   wire \add_x_19_4/n155 ;
   wire \add_x_19_4/n154 ;
   wire \add_x_19_4/n152 ;
   wire \add_x_19_4/n151 ;
   wire \add_x_19_4/n150 ;
   wire \add_x_19_4/n149 ;
   wire \add_x_19_4/n148 ;
   wire \add_x_19_4/n147 ;
   wire \add_x_19_4/n146 ;
   wire \add_x_19_4/n145 ;
   wire \add_x_19_4/n144 ;
   wire \add_x_19_4/n143 ;
   wire \add_x_19_4/n141 ;
   wire \add_x_19_4/n140 ;
   wire \add_x_19_4/n139 ;
   wire \add_x_19_4/n138 ;
   wire \add_x_19_4/n137 ;
   wire \add_x_19_4/n136 ;
   wire \add_x_19_4/n135 ;
   wire \add_x_19_4/n134 ;
   wire \add_x_19_4/n133 ;
   wire \add_x_19_4/n132 ;
   wire \add_x_19_4/n131 ;
   wire \add_x_19_4/n130 ;
   wire \add_x_19_4/n129 ;
   wire \add_x_19_4/n128 ;
   wire \add_x_19_4/n127 ;
   wire \add_x_19_4/n126 ;
   wire \add_x_19_4/n125 ;
   wire \add_x_19_4/n124 ;
   wire \add_x_19_4/n123 ;
   wire \add_x_19_4/n121 ;
   wire \add_x_19_4/n120 ;
   wire \add_x_19_4/n112 ;
   wire \add_x_19_4/n111 ;
   wire \add_x_19_4/n110 ;
   wire \add_x_19_4/n109 ;
   wire \add_x_19_4/n107 ;
   wire \add_x_19_4/n106 ;
   wire \add_x_19_4/n105 ;
   wire \add_x_19_4/n104 ;
   wire \add_x_19_4/n103 ;
   wire \add_x_19_4/n102 ;
   wire \add_x_19_4/n101 ;
   wire \add_x_19_4/n100 ;
   wire \add_x_19_4/n99 ;
   wire \add_x_19_4/n98 ;
   wire \add_x_19_4/n97 ;
   wire \add_x_19_4/n96 ;
   wire \add_x_19_4/n95 ;
   wire \add_x_19_4/n94 ;
   wire \add_x_19_4/n93 ;
   wire \add_x_19_4/n91 ;
   wire \add_x_19_4/n90 ;
   wire \add_x_19_4/n89 ;
   wire \add_x_19_4/n88 ;
   wire \add_x_19_4/n87 ;
   wire \add_x_19_4/n86 ;
   wire \add_x_19_4/n85 ;
   wire \add_x_19_4/n84 ;
   wire \add_x_19_4/n82 ;
   wire \add_x_19_4/n81 ;
   wire \add_x_19_4/n79 ;
   wire \add_x_19_4/n78 ;
   wire \add_x_19_4/n77 ;
   wire \add_x_19_4/n76 ;
   wire \add_x_19_4/n75 ;
   wire \add_x_19_4/n74 ;
   wire \add_x_19_4/n73 ;
   wire \add_x_19_4/n72 ;
   wire \add_x_19_4/n69 ;
   wire \add_x_19_4/n67 ;
   wire \add_x_19_4/n66 ;
   wire \add_x_19_4/n64 ;
   wire \add_x_19_4/n63 ;
   wire \add_x_19_4/n62 ;
   wire \add_x_19_4/n61 ;
   wire \add_x_19_4/n60 ;
   wire \add_x_19_4/n59 ;
   wire \add_x_19_4/n58 ;
   wire \add_x_19_4/n57 ;
   wire \add_x_19_4/n56 ;
   wire \add_x_19_4/n55 ;
   wire \add_x_19_4/n54 ;
   wire \add_x_19_4/n53 ;
   wire \add_x_19_4/n52 ;
   wire \add_x_19_4/n51 ;
   wire \add_x_19_4/n49 ;
   wire \add_x_19_4/n48 ;
   wire \add_x_19_4/n46 ;
   wire \add_x_19_4/n43 ;
   wire \add_x_19_4/n42 ;
   wire \add_x_19_4/n37 ;
   wire \add_x_19_4/n36 ;
   wire \add_x_19_4/n31 ;
   wire \add_x_19_4/n30 ;
   wire \add_x_19_4/n28 ;
   wire \add_x_19_4/n26 ;
   wire \add_x_19_4/n22 ;
   wire \add_x_19_4/n21 ;
   wire \add_x_19_4/n19 ;
   wire \add_x_19_4/n15 ;
   wire \add_x_19_4/n13 ;
   wire \add_x_19_4/n11 ;
   wire \add_x_19_4/n5 ;
   wire \add_x_19_4/n3 ;
   wire \add_x_19_2/n219 ;
   wire \add_x_19_2/n216 ;
   wire \add_x_19_2/n215 ;
   wire \add_x_19_2/n213 ;
   wire \add_x_19_2/n212 ;
   wire \add_x_19_2/n210 ;
   wire \add_x_19_2/n208 ;
   wire \add_x_19_2/n207 ;
   wire \add_x_19_2/n206 ;
   wire \add_x_19_2/n204 ;
   wire \add_x_19_2/n191 ;
   wire \add_x_19_2/n189 ;
   wire \add_x_19_2/n188 ;
   wire \add_x_19_2/n187 ;
   wire \add_x_19_2/n186 ;
   wire \add_x_19_2/n185 ;
   wire \add_x_19_2/n184 ;
   wire \add_x_19_2/n182 ;
   wire \add_x_19_2/n181 ;
   wire \add_x_19_2/n178 ;
   wire \add_x_19_2/n177 ;
   wire \add_x_19_2/n176 ;
   wire \add_x_19_2/n175 ;
   wire \add_x_19_2/n171 ;
   wire \add_x_19_2/n170 ;
   wire \add_x_19_2/n169 ;
   wire \add_x_19_2/n168 ;
   wire \add_x_19_2/n167 ;
   wire \add_x_19_2/n166 ;
   wire \add_x_19_2/n165 ;
   wire \add_x_19_2/n164 ;
   wire \add_x_19_2/n163 ;
   wire \add_x_19_2/n156 ;
   wire \add_x_19_2/n155 ;
   wire \add_x_19_2/n154 ;
   wire \add_x_19_2/n152 ;
   wire \add_x_19_2/n151 ;
   wire \add_x_19_2/n150 ;
   wire \add_x_19_2/n149 ;
   wire \add_x_19_2/n148 ;
   wire \add_x_19_2/n147 ;
   wire \add_x_19_2/n146 ;
   wire \add_x_19_2/n144 ;
   wire \add_x_19_2/n143 ;
   wire \add_x_19_2/n140 ;
   wire \add_x_19_2/n139 ;
   wire \add_x_19_2/n137 ;
   wire \add_x_19_2/n135 ;
   wire \add_x_19_2/n134 ;
   wire \add_x_19_2/n133 ;
   wire \add_x_19_2/n132 ;
   wire \add_x_19_2/n131 ;
   wire \add_x_19_2/n130 ;
   wire \add_x_19_2/n129 ;
   wire \add_x_19_2/n128 ;
   wire \add_x_19_2/n127 ;
   wire \add_x_19_2/n126 ;
   wire \add_x_19_2/n125 ;
   wire \add_x_19_2/n124 ;
   wire \add_x_19_2/n123 ;
   wire \add_x_19_2/n122 ;
   wire \add_x_19_2/n121 ;
   wire \add_x_19_2/n120 ;
   wire \add_x_19_2/n118 ;
   wire \add_x_19_2/n116 ;
   wire \add_x_19_2/n112 ;
   wire \add_x_19_2/n111 ;
   wire \add_x_19_2/n110 ;
   wire \add_x_19_2/n109 ;
   wire \add_x_19_2/n107 ;
   wire \add_x_19_2/n106 ;
   wire \add_x_19_2/n105 ;
   wire \add_x_19_2/n104 ;
   wire \add_x_19_2/n103 ;
   wire \add_x_19_2/n102 ;
   wire \add_x_19_2/n101 ;
   wire \add_x_19_2/n100 ;
   wire \add_x_19_2/n99 ;
   wire \add_x_19_2/n98 ;
   wire \add_x_19_2/n97 ;
   wire \add_x_19_2/n96 ;
   wire \add_x_19_2/n95 ;
   wire \add_x_19_2/n94 ;
   wire \add_x_19_2/n93 ;
   wire \add_x_19_2/n92 ;
   wire \add_x_19_2/n91 ;
   wire \add_x_19_2/n90 ;
   wire \add_x_19_2/n89 ;
   wire \add_x_19_2/n87 ;
   wire \add_x_19_2/n86 ;
   wire \add_x_19_2/n85 ;
   wire \add_x_19_2/n84 ;
   wire \add_x_19_2/n83 ;
   wire \add_x_19_2/n82 ;
   wire \add_x_19_2/n81 ;
   wire \add_x_19_2/n79 ;
   wire \add_x_19_2/n78 ;
   wire \add_x_19_2/n76 ;
   wire \add_x_19_2/n74 ;
   wire \add_x_19_2/n73 ;
   wire \add_x_19_2/n72 ;
   wire \add_x_19_2/n69 ;
   wire \add_x_19_2/n68 ;
   wire \add_x_19_2/n67 ;
   wire \add_x_19_2/n66 ;
   wire \add_x_19_2/n64 ;
   wire \add_x_19_2/n63 ;
   wire \add_x_19_2/n62 ;
   wire \add_x_19_2/n61 ;
   wire \add_x_19_2/n60 ;
   wire \add_x_19_2/n59 ;
   wire \add_x_19_2/n58 ;
   wire \add_x_19_2/n56 ;
   wire \add_x_19_2/n55 ;
   wire \add_x_19_2/n54 ;
   wire \add_x_19_2/n53 ;
   wire \add_x_19_2/n52 ;
   wire \add_x_19_2/n51 ;
   wire \add_x_19_2/n49 ;
   wire \add_x_19_2/n48 ;
   wire \add_x_19_2/n46 ;
   wire \add_x_19_2/n42 ;
   wire \add_x_19_2/n37 ;
   wire \add_x_19_2/n36 ;
   wire \add_x_19_2/n28 ;
   wire \add_x_19_2/n25 ;
   wire \add_x_19_2/n24 ;
   wire \add_x_19_2/n19 ;
   wire \add_x_19_2/n17 ;
   wire \add_x_19_2/n15 ;
   wire \add_x_19_1/n219 ;
   wire \add_x_19_1/n218 ;
   wire \add_x_19_1/n213 ;
   wire \add_x_19_1/n212 ;
   wire \add_x_19_1/n210 ;
   wire \add_x_19_1/n208 ;
   wire \add_x_19_1/n207 ;
   wire \add_x_19_1/n202 ;
   wire \add_x_19_1/n198 ;
   wire \add_x_19_1/n195 ;
   wire \add_x_19_1/n191 ;
   wire \add_x_19_1/n189 ;
   wire \add_x_19_1/n188 ;
   wire \add_x_19_1/n187 ;
   wire \add_x_19_1/n185 ;
   wire \add_x_19_1/n184 ;
   wire \add_x_19_1/n182 ;
   wire \add_x_19_1/n181 ;
   wire \add_x_19_1/n178 ;
   wire \add_x_19_1/n177 ;
   wire \add_x_19_1/n176 ;
   wire \add_x_19_1/n175 ;
   wire \add_x_19_1/n174 ;
   wire \add_x_19_1/n172 ;
   wire \add_x_19_1/n168 ;
   wire \add_x_19_1/n167 ;
   wire \add_x_19_1/n166 ;
   wire \add_x_19_1/n165 ;
   wire \add_x_19_1/n163 ;
   wire \add_x_19_1/n162 ;
   wire \add_x_19_1/n160 ;
   wire \add_x_19_1/n155 ;
   wire \add_x_19_1/n154 ;
   wire \add_x_19_1/n152 ;
   wire \add_x_19_1/n151 ;
   wire \add_x_19_1/n150 ;
   wire \add_x_19_1/n149 ;
   wire \add_x_19_1/n148 ;
   wire \add_x_19_1/n147 ;
   wire \add_x_19_1/n146 ;
   wire \add_x_19_1/n145 ;
   wire \add_x_19_1/n144 ;
   wire \add_x_19_1/n143 ;
   wire \add_x_19_1/n141 ;
   wire \add_x_19_1/n140 ;
   wire \add_x_19_1/n139 ;
   wire \add_x_19_1/n137 ;
   wire \add_x_19_1/n136 ;
   wire \add_x_19_1/n135 ;
   wire \add_x_19_1/n134 ;
   wire \add_x_19_1/n133 ;
   wire \add_x_19_1/n132 ;
   wire \add_x_19_1/n131 ;
   wire \add_x_19_1/n130 ;
   wire \add_x_19_1/n129 ;
   wire \add_x_19_1/n128 ;
   wire \add_x_19_1/n127 ;
   wire \add_x_19_1/n126 ;
   wire \add_x_19_1/n125 ;
   wire \add_x_19_1/n124 ;
   wire \add_x_19_1/n123 ;
   wire \add_x_19_1/n122 ;
   wire \add_x_19_1/n121 ;
   wire \add_x_19_1/n120 ;
   wire \add_x_19_1/n118 ;
   wire \add_x_19_1/n116 ;
   wire \add_x_19_1/n112 ;
   wire \add_x_19_1/n111 ;
   wire \add_x_19_1/n110 ;
   wire \add_x_19_1/n109 ;
   wire \add_x_19_1/n106 ;
   wire \add_x_19_1/n105 ;
   wire \add_x_19_1/n104 ;
   wire \add_x_19_1/n103 ;
   wire \add_x_19_1/n102 ;
   wire \add_x_19_1/n101 ;
   wire \add_x_19_1/n100 ;
   wire \add_x_19_1/n98 ;
   wire \add_x_19_1/n97 ;
   wire \add_x_19_1/n96 ;
   wire \add_x_19_1/n95 ;
   wire \add_x_19_1/n94 ;
   wire \add_x_19_1/n93 ;
   wire \add_x_19_1/n91 ;
   wire \add_x_19_1/n90 ;
   wire \add_x_19_1/n89 ;
   wire \add_x_19_1/n88 ;
   wire \add_x_19_1/n87 ;
   wire \add_x_19_1/n86 ;
   wire \add_x_19_1/n85 ;
   wire \add_x_19_1/n84 ;
   wire \add_x_19_1/n82 ;
   wire \add_x_19_1/n81 ;
   wire \add_x_19_1/n79 ;
   wire \add_x_19_1/n78 ;
   wire \add_x_19_1/n76 ;
   wire \add_x_19_1/n74 ;
   wire \add_x_19_1/n73 ;
   wire \add_x_19_1/n72 ;
   wire \add_x_19_1/n69 ;
   wire \add_x_19_1/n67 ;
   wire \add_x_19_1/n66 ;
   wire \add_x_19_1/n65 ;
   wire \add_x_19_1/n64 ;
   wire \add_x_19_1/n63 ;
   wire \add_x_19_1/n62 ;
   wire \add_x_19_1/n61 ;
   wire \add_x_19_1/n60 ;
   wire \add_x_19_1/n59 ;
   wire \add_x_19_1/n58 ;
   wire \add_x_19_1/n56 ;
   wire \add_x_19_1/n55 ;
   wire \add_x_19_1/n54 ;
   wire \add_x_19_1/n53 ;
   wire \add_x_19_1/n52 ;
   wire \add_x_19_1/n51 ;
   wire \add_x_19_1/n50 ;
   wire \add_x_19_1/n49 ;
   wire \add_x_19_1/n48 ;
   wire \add_x_19_1/n46 ;
   wire \add_x_19_1/n43 ;
   wire \add_x_19_1/n42 ;
   wire \add_x_19_1/n38 ;
   wire \add_x_19_1/n37 ;
   wire \add_x_19_1/n36 ;
   wire \add_x_19_1/n28 ;
   wire \add_x_19_1/n27 ;
   wire \add_x_19_1/n21 ;
   wire \add_x_19_1/n19 ;
   wire \add_x_19_1/n17 ;
   wire \add_x_19_1/n11 ;
   wire \add_x_19_1/n7 ;
   wire \add_x_19_1/n4 ;
   wire \add_x_19_1/n3 ;
   wire \add_x_19_3/n221 ;
   wire \add_x_19_3/n219 ;
   wire \add_x_19_3/n218 ;
   wire \add_x_19_3/n217 ;
   wire \add_x_19_3/n215 ;
   wire \add_x_19_3/n213 ;
   wire \add_x_19_3/n208 ;
   wire \add_x_19_3/n207 ;
   wire \add_x_19_3/n204 ;
   wire \add_x_19_3/n202 ;
   wire \add_x_19_3/n198 ;
   wire \add_x_19_3/n195 ;
   wire \add_x_19_3/n191 ;
   wire \add_x_19_3/n189 ;
   wire \add_x_19_3/n188 ;
   wire \add_x_19_3/n187 ;
   wire \add_x_19_3/n186 ;
   wire \add_x_19_3/n185 ;
   wire \add_x_19_3/n184 ;
   wire \add_x_19_3/n182 ;
   wire \add_x_19_3/n181 ;
   wire \add_x_19_3/n178 ;
   wire \add_x_19_3/n177 ;
   wire \add_x_19_3/n176 ;
   wire \add_x_19_3/n175 ;
   wire \add_x_19_3/n174 ;
   wire \add_x_19_3/n172 ;
   wire \add_x_19_3/n171 ;
   wire \add_x_19_3/n170 ;
   wire \add_x_19_3/n169 ;
   wire \add_x_19_3/n168 ;
   wire \add_x_19_3/n167 ;
   wire \add_x_19_3/n166 ;
   wire \add_x_19_3/n165 ;
   wire \add_x_19_3/n163 ;
   wire \add_x_19_3/n162 ;
   wire \add_x_19_3/n160 ;
   wire \add_x_19_3/n156 ;
   wire \add_x_19_3/n155 ;
   wire \add_x_19_3/n154 ;
   wire \add_x_19_3/n152 ;
   wire \add_x_19_3/n151 ;
   wire \add_x_19_3/n150 ;
   wire \add_x_19_3/n149 ;
   wire \add_x_19_3/n148 ;
   wire \add_x_19_3/n147 ;
   wire \add_x_19_3/n146 ;
   wire \add_x_19_3/n145 ;
   wire \add_x_19_3/n144 ;
   wire \add_x_19_3/n140 ;
   wire \add_x_19_3/n139 ;
   wire \add_x_19_3/n137 ;
   wire \add_x_19_3/n136 ;
   wire \add_x_19_3/n135 ;
   wire \add_x_19_3/n134 ;
   wire \add_x_19_3/n133 ;
   wire \add_x_19_3/n132 ;
   wire \add_x_19_3/n131 ;
   wire \add_x_19_3/n129 ;
   wire \add_x_19_3/n128 ;
   wire \add_x_19_3/n127 ;
   wire \add_x_19_3/n126 ;
   wire \add_x_19_3/n125 ;
   wire \add_x_19_3/n124 ;
   wire \add_x_19_3/n123 ;
   wire \add_x_19_3/n122 ;
   wire \add_x_19_3/n121 ;
   wire \add_x_19_3/n120 ;
   wire \add_x_19_3/n118 ;
   wire \add_x_19_3/n116 ;
   wire \add_x_19_3/n113 ;
   wire \add_x_19_3/n111 ;
   wire \add_x_19_3/n110 ;
   wire \add_x_19_3/n106 ;
   wire \add_x_19_3/n105 ;
   wire \add_x_19_3/n104 ;
   wire \add_x_19_3/n103 ;
   wire \add_x_19_3/n102 ;
   wire \add_x_19_3/n101 ;
   wire \add_x_19_3/n100 ;
   wire \add_x_19_3/n99 ;
   wire \add_x_19_3/n98 ;
   wire \add_x_19_3/n97 ;
   wire \add_x_19_3/n95 ;
   wire \add_x_19_3/n94 ;
   wire \add_x_19_3/n93 ;
   wire \add_x_19_3/n92 ;
   wire \add_x_19_3/n90 ;
   wire \add_x_19_3/n89 ;
   wire \add_x_19_3/n88 ;
   wire \add_x_19_3/n87 ;
   wire \add_x_19_3/n86 ;
   wire \add_x_19_3/n85 ;
   wire \add_x_19_3/n84 ;
   wire \add_x_19_3/n83 ;
   wire \add_x_19_3/n82 ;
   wire \add_x_19_3/n81 ;
   wire \add_x_19_3/n79 ;
   wire \add_x_19_3/n78 ;
   wire \add_x_19_3/n77 ;
   wire \add_x_19_3/n76 ;
   wire \add_x_19_3/n75 ;
   wire \add_x_19_3/n74 ;
   wire \add_x_19_3/n73 ;
   wire \add_x_19_3/n72 ;
   wire \add_x_19_3/n69 ;
   wire \add_x_19_3/n68 ;
   wire \add_x_19_3/n67 ;
   wire \add_x_19_3/n66 ;
   wire \add_x_19_3/n65 ;
   wire \add_x_19_3/n64 ;
   wire \add_x_19_3/n63 ;
   wire \add_x_19_3/n62 ;
   wire \add_x_19_3/n61 ;
   wire \add_x_19_3/n60 ;
   wire \add_x_19_3/n59 ;
   wire \add_x_19_3/n58 ;
   wire \add_x_19_3/n56 ;
   wire \add_x_19_3/n55 ;
   wire \add_x_19_3/n54 ;
   wire \add_x_19_3/n53 ;
   wire \add_x_19_3/n52 ;
   wire \add_x_19_3/n51 ;
   wire \add_x_19_3/n50 ;
   wire \add_x_19_3/n49 ;
   wire \add_x_19_3/n48 ;
   wire \add_x_19_3/n47 ;
   wire \add_x_19_3/n46 ;
   wire \add_x_19_3/n43 ;
   wire \add_x_19_3/n42 ;
   wire \add_x_19_3/n38 ;
   wire \add_x_19_3/n37 ;
   wire \add_x_19_3/n36 ;
   wire \add_x_19_3/n35 ;
   wire \add_x_19_3/n34 ;
   wire \add_x_19_3/n30 ;
   wire \add_x_19_3/n28 ;
   wire \add_x_19_3/n27 ;
   wire \add_x_19_3/n26 ;
   wire \add_x_19_3/n24 ;
   wire \add_x_19_3/n22 ;
   wire \add_x_19_3/n18 ;
   wire \add_x_19_3/n17 ;
   wire \add_x_19_3/n13 ;
   wire \add_x_19_3/n11 ;
   wire \add_x_19_3/n7 ;
   wire \add_x_19_3/n4 ;
   wire \add_x_19_5/n222 ;
   wire \add_x_19_5/n220 ;
   wire \add_x_19_5/n219 ;
   wire \add_x_19_5/n214 ;
   wire \add_x_19_5/n213 ;
   wire \add_x_19_5/n210 ;
   wire \add_x_19_5/n207 ;
   wire \add_x_19_5/n206 ;
   wire \add_x_19_5/n202 ;
   wire \add_x_19_5/n198 ;
   wire \add_x_19_5/n195 ;
   wire \add_x_19_5/n191 ;
   wire \add_x_19_5/n189 ;
   wire \add_x_19_5/n188 ;
   wire \add_x_19_5/n187 ;
   wire \add_x_19_5/n186 ;
   wire \add_x_19_5/n185 ;
   wire \add_x_19_5/n184 ;
   wire \add_x_19_5/n183 ;
   wire \add_x_19_5/n182 ;
   wire \add_x_19_5/n181 ;
   wire \add_x_19_5/n180 ;
   wire \add_x_19_5/n179 ;
   wire \add_x_19_5/n176 ;
   wire \add_x_19_5/n175 ;
   wire \add_x_19_5/n171 ;
   wire \add_x_19_5/n170 ;
   wire \add_x_19_5/n169 ;
   wire \add_x_19_5/n168 ;
   wire \add_x_19_5/n167 ;
   wire \add_x_19_5/n166 ;
   wire \add_x_19_5/n165 ;
   wire \add_x_19_5/n163 ;
   wire \add_x_19_5/n162 ;
   wire \add_x_19_5/n160 ;
   wire \add_x_19_5/n157 ;
   wire \add_x_19_5/n156 ;
   wire \add_x_19_5/n155 ;
   wire \add_x_19_5/n154 ;
   wire \add_x_19_5/n153 ;
   wire \add_x_19_5/n152 ;
   wire \add_x_19_5/n151 ;
   wire \add_x_19_5/n150 ;
   wire \add_x_19_5/n149 ;
   wire \add_x_19_5/n148 ;
   wire \add_x_19_5/n147 ;
   wire \add_x_19_5/n146 ;
   wire \add_x_19_5/n145 ;
   wire \add_x_19_5/n144 ;
   wire \add_x_19_5/n140 ;
   wire \add_x_19_5/n139 ;
   wire \add_x_19_5/n138 ;
   wire \add_x_19_5/n137 ;
   wire \add_x_19_5/n136 ;
   wire \add_x_19_5/n135 ;
   wire \add_x_19_5/n134 ;
   wire \add_x_19_5/n133 ;
   wire \add_x_19_5/n132 ;
   wire \add_x_19_5/n131 ;
   wire \add_x_19_5/n130 ;
   wire \add_x_19_5/n129 ;
   wire \add_x_19_5/n128 ;
   wire \add_x_19_5/n127 ;
   wire \add_x_19_5/n126 ;
   wire \add_x_19_5/n125 ;
   wire \add_x_19_5/n124 ;
   wire \add_x_19_5/n123 ;
   wire \add_x_19_5/n121 ;
   wire \add_x_19_5/n120 ;
   wire \add_x_19_5/n118 ;
   wire \add_x_19_5/n116 ;
   wire \add_x_19_5/n113 ;
   wire \add_x_19_5/n112 ;
   wire \add_x_19_5/n111 ;
   wire \add_x_19_5/n110 ;
   wire \add_x_19_5/n109 ;
   wire \add_x_19_5/n107 ;
   wire \add_x_19_5/n106 ;
   wire \add_x_19_5/n105 ;
   wire \add_x_19_5/n104 ;
   wire \add_x_19_5/n103 ;
   wire \add_x_19_5/n102 ;
   wire \add_x_19_5/n101 ;
   wire \add_x_19_5/n100 ;
   wire \add_x_19_5/n98 ;
   wire \add_x_19_5/n97 ;
   wire \add_x_19_5/n96 ;
   wire \add_x_19_5/n95 ;
   wire \add_x_19_5/n94 ;
   wire \add_x_19_5/n93 ;
   wire \add_x_19_5/n92 ;
   wire \add_x_19_5/n91 ;
   wire \add_x_19_5/n90 ;
   wire \add_x_19_5/n89 ;
   wire \add_x_19_5/n88 ;
   wire \add_x_19_5/n87 ;
   wire \add_x_19_5/n86 ;
   wire \add_x_19_5/n85 ;
   wire \add_x_19_5/n84 ;
   wire \add_x_19_5/n83 ;
   wire \add_x_19_5/n82 ;
   wire \add_x_19_5/n81 ;
   wire \add_x_19_5/n79 ;
   wire \add_x_19_5/n78 ;
   wire \add_x_19_5/n76 ;
   wire \add_x_19_5/n74 ;
   wire \add_x_19_5/n73 ;
   wire \add_x_19_5/n72 ;
   wire \add_x_19_5/n69 ;
   wire \add_x_19_5/n68 ;
   wire \add_x_19_5/n67 ;
   wire \add_x_19_5/n66 ;
   wire \add_x_19_5/n65 ;
   wire \add_x_19_5/n64 ;
   wire \add_x_19_5/n63 ;
   wire \add_x_19_5/n62 ;
   wire \add_x_19_5/n61 ;
   wire \add_x_19_5/n60 ;
   wire \add_x_19_5/n59 ;
   wire \add_x_19_5/n58 ;
   wire \add_x_19_5/n56 ;
   wire \add_x_19_5/n55 ;
   wire \add_x_19_5/n53 ;
   wire \add_x_19_5/n52 ;
   wire \add_x_19_5/n51 ;
   wire \add_x_19_5/n50 ;
   wire \add_x_19_5/n49 ;
   wire \add_x_19_5/n48 ;
   wire \add_x_19_5/n46 ;
   wire \add_x_19_5/n43 ;
   wire \add_x_19_5/n42 ;
   wire \add_x_19_5/n37 ;
   wire \add_x_19_5/n36 ;
   wire \add_x_19_5/n31 ;
   wire \add_x_19_5/n29 ;
   wire \add_x_19_5/n28 ;
   wire \add_x_19_5/n23 ;
   wire \add_x_19_5/n22 ;
   wire \add_x_19_5/n19 ;
   wire \add_x_19_5/n16 ;
   wire \add_x_19_5/n15 ;
   wire \add_x_19_5/n11 ;
   wire \add_x_19_5/n7 ;
   wire \add_x_19_5/n4 ;
   wire \add_x_19_0/n219 ;
   wire \add_x_19_0/n215 ;
   wire \add_x_19_0/n213 ;
   wire \add_x_19_0/n210 ;
   wire \add_x_19_0/n208 ;
   wire \add_x_19_0/n207 ;
   wire \add_x_19_0/n206 ;
   wire \add_x_19_0/n204 ;
   wire \add_x_19_0/n202 ;
   wire \add_x_19_0/n198 ;
   wire \add_x_19_0/n195 ;
   wire \add_x_19_0/n191 ;
   wire \add_x_19_0/n189 ;
   wire \add_x_19_0/n188 ;
   wire \add_x_19_0/n187 ;
   wire \add_x_19_0/n186 ;
   wire \add_x_19_0/n185 ;
   wire \add_x_19_0/n184 ;
   wire \add_x_19_0/n182 ;
   wire \add_x_19_0/n181 ;
   wire \add_x_19_0/n178 ;
   wire \add_x_19_0/n177 ;
   wire \add_x_19_0/n176 ;
   wire \add_x_19_0/n175 ;
   wire \add_x_19_0/n171 ;
   wire \add_x_19_0/n170 ;
   wire \add_x_19_0/n169 ;
   wire \add_x_19_0/n168 ;
   wire \add_x_19_0/n167 ;
   wire \add_x_19_0/n166 ;
   wire \add_x_19_0/n165 ;
   wire \add_x_19_0/n163 ;
   wire \add_x_19_0/n162 ;
   wire \add_x_19_0/n156 ;
   wire \add_x_19_0/n155 ;
   wire \add_x_19_0/n154 ;
   wire \add_x_19_0/n152 ;
   wire \add_x_19_0/n151 ;
   wire \add_x_19_0/n150 ;
   wire \add_x_19_0/n149 ;
   wire \add_x_19_0/n148 ;
   wire \add_x_19_0/n147 ;
   wire \add_x_19_0/n146 ;
   wire \add_x_19_0/n145 ;
   wire \add_x_19_0/n144 ;
   wire \add_x_19_0/n140 ;
   wire \add_x_19_0/n139 ;
   wire \add_x_19_0/n137 ;
   wire \add_x_19_0/n136 ;
   wire \add_x_19_0/n135 ;
   wire \add_x_19_0/n133 ;
   wire \add_x_19_0/n132 ;
   wire \add_x_19_0/n131 ;
   wire \add_x_19_0/n130 ;
   wire \add_x_19_0/n129 ;
   wire \add_x_19_0/n128 ;
   wire \add_x_19_0/n127 ;
   wire \add_x_19_0/n126 ;
   wire \add_x_19_0/n125 ;
   wire \add_x_19_0/n124 ;
   wire \add_x_19_0/n123 ;
   wire \add_x_19_0/n122 ;
   wire \add_x_19_0/n121 ;
   wire \add_x_19_0/n120 ;
   wire \add_x_19_0/n118 ;
   wire \add_x_19_0/n112 ;
   wire \add_x_19_0/n111 ;
   wire \add_x_19_0/n110 ;
   wire \add_x_19_0/n109 ;
   wire \add_x_19_0/n107 ;
   wire \add_x_19_0/n106 ;
   wire \add_x_19_0/n105 ;
   wire \add_x_19_0/n104 ;
   wire \add_x_19_0/n103 ;
   wire \add_x_19_0/n102 ;
   wire \add_x_19_0/n101 ;
   wire \add_x_19_0/n100 ;
   wire \add_x_19_0/n99 ;
   wire \add_x_19_0/n98 ;
   wire \add_x_19_0/n97 ;
   wire \add_x_19_0/n95 ;
   wire \add_x_19_0/n94 ;
   wire \add_x_19_0/n93 ;
   wire \add_x_19_0/n90 ;
   wire \add_x_19_0/n89 ;
   wire \add_x_19_0/n88 ;
   wire \add_x_19_0/n87 ;
   wire \add_x_19_0/n86 ;
   wire \add_x_19_0/n85 ;
   wire \add_x_19_0/n84 ;
   wire \add_x_19_0/n82 ;
   wire \add_x_19_0/n81 ;
   wire \add_x_19_0/n79 ;
   wire \add_x_19_0/n78 ;
   wire \add_x_19_0/n76 ;
   wire \add_x_19_0/n74 ;
   wire \add_x_19_0/n73 ;
   wire \add_x_19_0/n72 ;
   wire \add_x_19_0/n69 ;
   wire \add_x_19_0/n68 ;
   wire \add_x_19_0/n67 ;
   wire \add_x_19_0/n66 ;
   wire \add_x_19_0/n65 ;
   wire \add_x_19_0/n64 ;
   wire \add_x_19_0/n63 ;
   wire \add_x_19_0/n62 ;
   wire \add_x_19_0/n61 ;
   wire \add_x_19_0/n60 ;
   wire \add_x_19_0/n59 ;
   wire \add_x_19_0/n58 ;
   wire \add_x_19_0/n56 ;
   wire \add_x_19_0/n55 ;
   wire \add_x_19_0/n54 ;
   wire \add_x_19_0/n53 ;
   wire \add_x_19_0/n52 ;
   wire \add_x_19_0/n51 ;
   wire \add_x_19_0/n50 ;
   wire \add_x_19_0/n49 ;
   wire \add_x_19_0/n48 ;
   wire \add_x_19_0/n47 ;
   wire \add_x_19_0/n46 ;
   wire \add_x_19_0/n45 ;
   wire \add_x_19_0/n44 ;
   wire \add_x_19_0/n43 ;
   wire \add_x_19_0/n42 ;
   wire \add_x_19_0/n38 ;
   wire \add_x_19_0/n37 ;
   wire \add_x_19_0/n36 ;
   wire \add_x_19_0/n34 ;
   wire \add_x_19_0/n28 ;
   wire \add_x_19_0/n24 ;
   wire \add_x_19_0/n22 ;
   wire \add_x_19_0/n19 ;
   wire \add_x_19_0/n17 ;
   wire \add_x_19_0/n15 ;
   wire \add_x_19_0/n13 ;
   wire \add_x_19_0/n11 ;
   wire \add_x_19_0/n7 ;
   wire \add_x_19_0/n4 ;
   wire \add_x_19_0/n1 ;
   wire \DP_OP_159_297_3515/n1138 ;
   wire \DP_OP_159_297_3515/n1133 ;
   wire \DP_OP_159_297_3515/n1128 ;
   wire \DP_OP_159_297_3515/n1074 ;
   wire \DP_OP_159_297_3515/n1069 ;
   wire \DP_OP_159_297_3515/n1064 ;
   wire \DP_OP_159_297_3515/n1063 ;
   wire \DP_OP_159_297_3515/n1057 ;
   wire \DP_OP_159_297_3515/n1052 ;
   wire \DP_OP_159_297_3515/n1051 ;
   wire \DP_OP_159_297_3515/n1044 ;
   wire \DP_OP_159_297_3515/n1039 ;
   wire \DP_OP_159_297_3515/n1031 ;
   wire \DP_OP_159_297_3515/n1026 ;
   wire \DP_OP_159_297_3515/n1025 ;
   wire \DP_OP_159_297_3515/n1024 ;
   wire \DP_OP_159_297_3515/n1018 ;
   wire \DP_OP_159_297_3515/n1017 ;
   wire \DP_OP_159_297_3515/n1012 ;
   wire \DP_OP_159_297_3515/n1011 ;
   wire \DP_OP_159_297_3515/n1010 ;
   wire \DP_OP_159_297_3515/n1004 ;
   wire \DP_OP_159_297_3515/n1003 ;
   wire \DP_OP_159_297_3515/n999 ;
   wire \DP_OP_159_297_3515/n998 ;
   wire \DP_OP_159_297_3515/n997 ;
   wire \DP_OP_159_297_3515/n996 ;
   wire \DP_OP_159_297_3515/n991 ;
   wire \DP_OP_159_297_3515/n990 ;
   wire \DP_OP_159_297_3515/n989 ;
   wire \DP_OP_159_297_3515/n976 ;
   wire \DP_OP_159_297_3515/n971 ;
   wire \DP_OP_159_297_3515/n964 ;
   wire \DP_OP_159_297_3515/n963 ;
   wire \DP_OP_159_297_3515/n959 ;
   wire \DP_OP_159_297_3515/n957 ;
   wire \DP_OP_159_297_3515/n956 ;
   wire \DP_OP_159_297_3515/n955 ;
   wire \DP_OP_159_297_3515/n950 ;
   wire \DP_OP_159_297_3515/n949 ;
   wire \DP_OP_159_297_3515/n948 ;
   wire \DP_OP_159_297_3515/n944 ;
   wire \DP_OP_159_297_3515/n943 ;
   wire \DP_OP_159_297_3515/n936 ;
   wire \DP_OP_159_297_3515/n935 ;
   wire \DP_OP_159_297_3515/n934 ;
   wire \DP_OP_159_297_3515/n931 ;
   wire \DP_OP_159_297_3515/n930 ;
   wire \DP_OP_159_297_3515/n928 ;
   wire \DP_OP_159_297_3515/n927 ;
   wire \DP_OP_159_297_3515/n921 ;
   wire \DP_OP_159_297_3515/n920 ;
   wire \DP_OP_159_297_3515/n916 ;
   wire \DP_OP_159_297_3515/n915 ;
   wire \DP_OP_159_297_3515/n914 ;
   wire \DP_OP_159_297_3515/n913 ;
   wire \DP_OP_159_297_3515/n908 ;
   wire \DP_OP_159_297_3515/n907 ;
   wire \DP_OP_159_297_3515/n906 ;
   wire \DP_OP_159_297_3515/n902 ;
   wire \DP_OP_159_297_3515/n894 ;
   wire \DP_OP_159_297_3515/n893 ;
   wire \DP_OP_159_297_3515/n892 ;
   wire \DP_OP_159_297_3515/n887 ;
   wire \DP_OP_159_297_3515/n886 ;
   wire \DP_OP_159_297_3515/n885 ;
   wire \DP_OP_159_297_3515/n880 ;
   wire \DP_OP_159_297_3515/n879 ;
   wire \DP_OP_159_297_3515/n878 ;
   wire \DP_OP_159_297_3515/n877 ;
   wire \DP_OP_159_297_3515/n876 ;
   wire \DP_OP_159_297_3515/n875 ;
   wire \DP_OP_159_297_3515/n873 ;
   wire \DP_OP_159_297_3515/n871 ;
   wire \DP_OP_159_297_3515/n870 ;
   wire \DP_OP_159_297_3515/n869 ;
   wire \DP_OP_159_297_3515/n867 ;
   wire \DP_OP_159_297_3515/n862 ;
   wire \DP_OP_159_297_3515/n852 ;
   wire \DP_OP_159_297_3515/n815 ;
   wire \DP_OP_159_297_3515/n778 ;
   wire \DP_OP_159_297_3515/n776 ;
   wire \DP_OP_159_297_3515/n774 ;
   wire \DP_OP_159_297_3515/n768 ;
   wire \DP_OP_159_297_3515/n766 ;
   wire \DP_OP_159_297_3515/n764 ;
   wire \DP_OP_159_297_3515/n758 ;
   wire \DP_OP_159_297_3515/n742 ;
   wire \DP_OP_159_297_3515/n740 ;
   wire \DP_OP_159_297_3515/n737 ;
   wire \DP_OP_159_297_3515/n730 ;
   wire \DP_OP_159_297_3515/n728 ;
   wire \DP_OP_159_297_3515/n726 ;
   wire \DP_OP_159_297_3515/n723 ;
   wire \DP_OP_159_297_3515/n714 ;
   wire \DP_OP_159_297_3515/n712 ;
   wire \DP_OP_159_297_3515/n705 ;
   wire \DP_OP_159_297_3515/n694 ;
   wire \DP_OP_159_297_3515/n692 ;
   wire \DP_OP_159_297_3515/n690 ;
   wire \DP_OP_159_297_3515/n688 ;
   wire \DP_OP_159_297_3515/n685 ;
   wire \DP_OP_159_297_3515/n674 ;
   wire \DP_OP_159_297_3515/n672 ;
   wire \DP_OP_159_297_3515/n650 ;
   wire \DP_OP_159_297_3515/n648 ;
   wire \DP_OP_159_297_3515/n646 ;
   wire \DP_OP_159_297_3515/n638 ;
   wire \DP_OP_159_297_3515/n625 ;
   wire \DP_OP_159_297_3515/n623 ;
   wire \DP_OP_159_297_3515/n610 ;
   wire \DP_OP_159_297_3515/n593 ;
   wire \DP_OP_159_297_3515/n591 ;
   wire \DP_OP_159_297_3515/n589 ;
   wire \DP_OP_159_297_3515/n587 ;
   wire \DP_OP_159_297_3515/n160 ;
   wire \DP_OP_159_297_3515/n1 ;
   wire \DP_OP_158_296_6262/n2060 ;
   wire \DP_OP_158_296_6262/n2054 ;
   wire \DP_OP_158_296_6262/n2051 ;
   wire \DP_OP_158_296_6262/n2048 ;
   wire \DP_OP_158_296_6262/n2034 ;
   wire \DP_OP_158_296_6262/n2020 ;
   wire \DP_OP_158_296_6262/n2015 ;
   wire \DP_OP_158_296_6262/n2011 ;
   wire \DP_OP_158_296_6262/n2010 ;
   wire \DP_OP_158_296_6262/n2004 ;
   wire \DP_OP_158_296_6262/n1999 ;
   wire \DP_OP_158_296_6262/n1998 ;
   wire \DP_OP_158_296_6262/n1991 ;
   wire \DP_OP_158_296_6262/n1987 ;
   wire \DP_OP_158_296_6262/n1978 ;
   wire \DP_OP_158_296_6262/n1973 ;
   wire \DP_OP_158_296_6262/n1972 ;
   wire \DP_OP_158_296_6262/n1971 ;
   wire \DP_OP_158_296_6262/n1966 ;
   wire \DP_OP_158_296_6262/n1965 ;
   wire \DP_OP_158_296_6262/n1964 ;
   wire \DP_OP_158_296_6262/n1959 ;
   wire \DP_OP_158_296_6262/n1958 ;
   wire \DP_OP_158_296_6262/n1957 ;
   wire \DP_OP_158_296_6262/n1952 ;
   wire \DP_OP_158_296_6262/n1951 ;
   wire \DP_OP_158_296_6262/n1950 ;
   wire \DP_OP_158_296_6262/n1946 ;
   wire \DP_OP_158_296_6262/n1945 ;
   wire \DP_OP_158_296_6262/n1944 ;
   wire \DP_OP_158_296_6262/n1943 ;
   wire \DP_OP_158_296_6262/n1938 ;
   wire \DP_OP_158_296_6262/n1937 ;
   wire \DP_OP_158_296_6262/n1936 ;
   wire \DP_OP_158_296_6262/n1918 ;
   wire \DP_OP_158_296_6262/n1917 ;
   wire \DP_OP_158_296_6262/n1916 ;
   wire \DP_OP_158_296_6262/n1911 ;
   wire \DP_OP_158_296_6262/n1910 ;
   wire \DP_OP_158_296_6262/n1909 ;
   wire \DP_OP_158_296_6262/n1904 ;
   wire \DP_OP_158_296_6262/n1903 ;
   wire \DP_OP_158_296_6262/n1897 ;
   wire \DP_OP_158_296_6262/n1896 ;
   wire \DP_OP_158_296_6262/n1895 ;
   wire \DP_OP_158_296_6262/n1890 ;
   wire \DP_OP_158_296_6262/n1881 ;
   wire \DP_OP_158_296_6262/n1877 ;
   wire \DP_OP_158_296_6262/n1875 ;
   wire \DP_OP_158_296_6262/n1874 ;
   wire \DP_OP_158_296_6262/n1869 ;
   wire \DP_OP_158_296_6262/n1863 ;
   wire \DP_OP_158_296_6262/n1862 ;
   wire \DP_OP_158_296_6262/n1855 ;
   wire \DP_OP_158_296_6262/n1854 ;
   wire \DP_OP_158_296_6262/n1849 ;
   wire \DP_OP_158_296_6262/n1848 ;
   wire \DP_OP_158_296_6262/n1847 ;
   wire \DP_OP_158_296_6262/n1837 ;
   wire \DP_OP_158_296_6262/n1834 ;
   wire \DP_OP_158_296_6262/n1833 ;
   wire \DP_OP_158_296_6262/n1830 ;
   wire \DP_OP_158_296_6262/n1829 ;
   wire \DP_OP_158_296_6262/n1828 ;
   wire \DP_OP_158_296_6262/n1827 ;
   wire \DP_OP_158_296_6262/n1826 ;
   wire \DP_OP_158_296_6262/n1792 ;
   wire \DP_OP_158_296_6262/n1791 ;
   wire \DP_OP_158_296_6262/n855 ;
   wire \DP_OP_158_296_6262/n841 ;
   wire \DP_OP_158_296_6262/n838 ;
   wire \DP_OP_158_296_6262/n833 ;
   wire \DP_OP_158_296_6262/n829 ;
   wire \DP_OP_158_296_6262/n375 ;
   wire \DP_OP_158_296_6262/n373 ;
   wire \DP_OP_158_296_6262/n371 ;
   wire \DP_OP_158_296_6262/n365 ;
   wire \DP_OP_158_296_6262/n349 ;
   wire \DP_OP_158_296_6262/n347 ;
   wire \DP_OP_158_296_6262/n329 ;
   wire \DP_OP_158_296_6262/n322 ;
   wire \DP_OP_158_296_6262/n320 ;
   wire \DP_OP_158_296_6262/n318 ;
   wire \DP_OP_158_296_6262/n315 ;
   wire \DP_OP_158_296_6262/n306 ;
   wire \DP_OP_158_296_6262/n304 ;
   wire \DP_OP_158_296_6262/n297 ;
   wire \DP_OP_158_296_6262/n286 ;
   wire \DP_OP_158_296_6262/n284 ;
   wire \DP_OP_158_296_6262/n282 ;
   wire \DP_OP_158_296_6262/n280 ;
   wire \DP_OP_158_296_6262/n277 ;
   wire \DP_OP_158_296_6262/n266 ;
   wire \DP_OP_158_296_6262/n264 ;
   wire \DP_OP_158_296_6262/n255 ;
   wire \DP_OP_158_296_6262/n242 ;
   wire \DP_OP_158_296_6262/n240 ;
   wire \DP_OP_158_296_6262/n238 ;
   wire \DP_OP_158_296_6262/n230 ;
   wire \DP_OP_158_296_6262/n217 ;
   wire \DP_OP_158_296_6262/n215 ;
   wire \DP_OP_158_296_6262/n202 ;
   wire \DP_OP_158_296_6262/n185 ;
   wire \DP_OP_158_296_6262/n183 ;
   wire \DP_OP_158_296_6262/n181 ;
   wire \DP_OP_158_296_6262/n179 ;
   wire \DP_OP_158_296_6262/n174 ;
   wire \DP_OP_158_296_6262/n161 ;
   wire \DP_OP_158_296_6262/n159 ;
   wire \DP_OP_158_296_6262/n148 ;
   wire \DP_OP_158_296_6262/n133 ;
   wire \DP_OP_158_296_6262/n131 ;
   wire \DP_OP_158_296_6262/n129 ;
   wire \DP_OP_158_296_6262/n119 ;
   wire \DP_OP_158_296_6262/n104 ;
   wire \DP_OP_158_296_6262/n102 ;
   wire \DP_OP_158_296_6262/n87 ;
   wire \DP_OP_158_296_6262/n68 ;
   wire \DP_OP_158_296_6262/n66 ;
   wire \DP_OP_158_296_6262/n64 ;
   wire \DP_OP_158_296_6262/n62 ;
   wire \DP_OP_158_296_6262/n54 ;
   wire \DP_OP_158_296_6262/n39 ;
   wire \DP_OP_158_296_6262/n37 ;
   wire \DP_OP_158_296_6262/n18 ;
   wire \DP_OP_158_296_6262/n5 ;
   wire \DP_OP_158_296_6262/n3 ;
   wire \add_x_22_4/n121 ;
   wire \add_x_22_4/n119 ;
   wire \add_x_22_4/n118 ;
   wire \add_x_22_4/n117 ;
   wire \add_x_22_4/n115 ;
   wire \add_x_22_4/n112 ;
   wire \add_x_22_4/n111 ;
   wire \add_x_22_4/n110 ;
   wire \add_x_22_4/n109 ;
   wire \add_x_22_4/n106 ;
   wire \add_x_22_4/n105 ;
   wire \add_x_22_4/n103 ;
   wire \add_x_22_4/n102 ;
   wire \add_x_22_4/n101 ;
   wire \add_x_22_4/n99 ;
   wire \add_x_22_4/n98 ;
   wire \add_x_22_4/n94 ;
   wire \add_x_22_4/n93 ;
   wire \add_x_22_4/n92 ;
   wire \add_x_22_4/n90 ;
   wire \add_x_22_4/n87 ;
   wire \add_x_22_4/n85 ;
   wire \add_x_22_4/n84 ;
   wire \add_x_22_4/n81 ;
   wire \add_x_22_4/n80 ;
   wire \add_x_22_4/n78 ;
   wire \add_x_22_4/n77 ;
   wire \add_x_22_4/n76 ;
   wire \add_x_22_4/n75 ;
   wire \add_x_22_4/n74 ;
   wire \add_x_22_4/n71 ;
   wire \add_x_22_4/n69 ;
   wire \add_x_22_4/n68 ;
   wire \add_x_22_4/n67 ;
   wire \add_x_22_4/n65 ;
   wire \add_x_22_4/n64 ;
   wire \add_x_22_4/n59 ;
   wire \add_x_22_4/n58 ;
   wire \add_x_22_4/n57 ;
   wire \add_x_22_4/n54 ;
   wire \add_x_22_4/n51 ;
   wire \add_x_22_4/n50 ;
   wire \add_x_22_4/n47 ;
   wire \add_x_22_4/n46 ;
   wire \add_x_22_4/n44 ;
   wire \add_x_22_4/n43 ;
   wire \add_x_22_4/n42 ;
   wire \add_x_22_4/n41 ;
   wire \add_x_22_4/n35 ;
   wire \add_x_22_4/n34 ;
   wire \add_x_22_4/n33 ;
   wire \add_x_22_4/n30 ;
   wire \add_x_22_4/n28 ;
   wire \add_x_22_4/n27 ;
   wire \add_x_22_4/n26 ;
   wire \add_x_22_4/n24 ;
   wire \add_x_22_4/n23 ;
   wire \add_x_22_4/n20 ;
   wire \add_x_22_4/n17 ;
   wire \add_x_22_4/n16 ;
   wire \add_x_22_4/n15 ;
   wire \add_x_22_4/n10 ;
   wire \add_x_22_4/n9 ;
   wire \add_x_22_4/n8 ;
   wire \add_x_22_4/n7 ;
   wire \add_x_22_4/n2 ;
   wire \add_x_22_4/n1 ;
   wire \add_x_22_1/n121 ;
   wire \add_x_22_1/n119 ;
   wire \add_x_22_1/n118 ;
   wire \add_x_22_1/n117 ;
   wire \add_x_22_1/n115 ;
   wire \add_x_22_1/n114 ;
   wire \add_x_22_1/n112 ;
   wire \add_x_22_1/n111 ;
   wire \add_x_22_1/n110 ;
   wire \add_x_22_1/n109 ;
   wire \add_x_22_1/n103 ;
   wire \add_x_22_1/n102 ;
   wire \add_x_22_1/n99 ;
   wire \add_x_22_1/n98 ;
   wire \add_x_22_1/n96 ;
   wire \add_x_22_1/n95 ;
   wire \add_x_22_1/n94 ;
   wire \add_x_22_1/n93 ;
   wire \add_x_22_1/n92 ;
   wire \add_x_22_1/n90 ;
   wire \add_x_22_1/n89 ;
   wire \add_x_22_1/n87 ;
   wire \add_x_22_1/n85 ;
   wire \add_x_22_1/n84 ;
   wire \add_x_22_1/n78 ;
   wire \add_x_22_1/n77 ;
   wire \add_x_22_1/n76 ;
   wire \add_x_22_1/n75 ;
   wire \add_x_22_1/n74 ;
   wire \add_x_22_1/n72 ;
   wire \add_x_22_1/n71 ;
   wire \add_x_22_1/n69 ;
   wire \add_x_22_1/n68 ;
   wire \add_x_22_1/n67 ;
   wire \add_x_22_1/n65 ;
   wire \add_x_22_1/n64 ;
   wire \add_x_22_1/n59 ;
   wire \add_x_22_1/n58 ;
   wire \add_x_22_1/n57 ;
   wire \add_x_22_1/n54 ;
   wire \add_x_22_1/n53 ;
   wire \add_x_22_1/n51 ;
   wire \add_x_22_1/n50 ;
   wire \add_x_22_1/n47 ;
   wire \add_x_22_1/n44 ;
   wire \add_x_22_1/n43 ;
   wire \add_x_22_1/n42 ;
   wire \add_x_22_1/n41 ;
   wire \add_x_22_1/n38 ;
   wire \add_x_22_1/n35 ;
   wire \add_x_22_1/n34 ;
   wire \add_x_22_1/n31 ;
   wire \add_x_22_1/n30 ;
   wire \add_x_22_1/n28 ;
   wire \add_x_22_1/n27 ;
   wire \add_x_22_1/n26 ;
   wire \add_x_22_1/n24 ;
   wire \add_x_22_1/n23 ;
   wire \add_x_22_1/n20 ;
   wire \add_x_22_1/n17 ;
   wire \add_x_22_1/n16 ;
   wire \add_x_22_1/n15 ;
   wire \add_x_22_1/n10 ;
   wire \add_x_22_1/n9 ;
   wire \add_x_22_1/n8 ;
   wire \add_x_22_1/n7 ;
   wire \add_x_22_1/n5 ;
   wire \add_x_22_1/n4 ;
   wire \add_x_22_1/n3 ;
   wire \add_x_22_1/n2 ;
   wire \add_x_22_1/n1 ;
   wire \add_x_22_5/n121 ;
   wire \add_x_22_5/n119 ;
   wire \add_x_22_5/n118 ;
   wire \add_x_22_5/n117 ;
   wire \add_x_22_5/n115 ;
   wire \add_x_22_5/n114 ;
   wire \add_x_22_5/n112 ;
   wire \add_x_22_5/n111 ;
   wire \add_x_22_5/n110 ;
   wire \add_x_22_5/n109 ;
   wire \add_x_22_5/n106 ;
   wire \add_x_22_5/n103 ;
   wire \add_x_22_5/n102 ;
   wire \add_x_22_5/n101 ;
   wire \add_x_22_5/n99 ;
   wire \add_x_22_5/n94 ;
   wire \add_x_22_5/n93 ;
   wire \add_x_22_5/n92 ;
   wire \add_x_22_5/n90 ;
   wire \add_x_22_5/n89 ;
   wire \add_x_22_5/n87 ;
   wire \add_x_22_5/n85 ;
   wire \add_x_22_5/n84 ;
   wire \add_x_22_5/n81 ;
   wire \add_x_22_5/n80 ;
   wire \add_x_22_5/n78 ;
   wire \add_x_22_5/n77 ;
   wire \add_x_22_5/n76 ;
   wire \add_x_22_5/n75 ;
   wire \add_x_22_5/n74 ;
   wire \add_x_22_5/n72 ;
   wire \add_x_22_5/n71 ;
   wire \add_x_22_5/n69 ;
   wire \add_x_22_5/n68 ;
   wire \add_x_22_5/n67 ;
   wire \add_x_22_5/n59 ;
   wire \add_x_22_5/n58 ;
   wire \add_x_22_5/n57 ;
   wire \add_x_22_5/n54 ;
   wire \add_x_22_5/n53 ;
   wire \add_x_22_5/n51 ;
   wire \add_x_22_5/n50 ;
   wire \add_x_22_5/n47 ;
   wire \add_x_22_5/n44 ;
   wire \add_x_22_5/n43 ;
   wire \add_x_22_5/n42 ;
   wire \add_x_22_5/n41 ;
   wire \add_x_22_5/n35 ;
   wire \add_x_22_5/n34 ;
   wire \add_x_22_5/n33 ;
   wire \add_x_22_5/n31 ;
   wire \add_x_22_5/n26 ;
   wire \add_x_22_5/n24 ;
   wire \add_x_22_5/n23 ;
   wire \add_x_22_5/n20 ;
   wire \add_x_22_5/n17 ;
   wire \add_x_22_5/n16 ;
   wire \add_x_22_5/n15 ;
   wire \add_x_22_5/n13 ;
   wire \add_x_22_5/n10 ;
   wire \add_x_22_5/n9 ;
   wire \add_x_22_5/n8 ;
   wire \add_x_22_5/n5 ;
   wire \add_x_22_5/n4 ;
   wire \add_x_22_5/n3 ;
   wire \add_x_22_5/n2 ;
   wire \add_x_22_5/n1 ;
   wire \add_x_22_3/n119 ;
   wire \add_x_22_3/n118 ;
   wire \add_x_22_3/n115 ;
   wire \add_x_22_3/n114 ;
   wire \add_x_22_3/n112 ;
   wire \add_x_22_3/n111 ;
   wire \add_x_22_3/n110 ;
   wire \add_x_22_3/n109 ;
   wire \add_x_22_3/n106 ;
   wire \add_x_22_3/n105 ;
   wire \add_x_22_3/n103 ;
   wire \add_x_22_3/n102 ;
   wire \add_x_22_3/n101 ;
   wire \add_x_22_3/n98 ;
   wire \add_x_22_3/n94 ;
   wire \add_x_22_3/n93 ;
   wire \add_x_22_3/n92 ;
   wire \add_x_22_3/n90 ;
   wire \add_x_22_3/n89 ;
   wire \add_x_22_3/n87 ;
   wire \add_x_22_3/n85 ;
   wire \add_x_22_3/n84 ;
   wire \add_x_22_3/n81 ;
   wire \add_x_22_3/n80 ;
   wire \add_x_22_3/n78 ;
   wire \add_x_22_3/n77 ;
   wire \add_x_22_3/n76 ;
   wire \add_x_22_3/n75 ;
   wire \add_x_22_3/n72 ;
   wire \add_x_22_3/n71 ;
   wire \add_x_22_3/n69 ;
   wire \add_x_22_3/n68 ;
   wire \add_x_22_3/n59 ;
   wire \add_x_22_3/n58 ;
   wire \add_x_22_3/n57 ;
   wire \add_x_22_3/n54 ;
   wire \add_x_22_3/n51 ;
   wire \add_x_22_3/n50 ;
   wire \add_x_22_3/n47 ;
   wire \add_x_22_3/n44 ;
   wire \add_x_22_3/n43 ;
   wire \add_x_22_3/n42 ;
   wire \add_x_22_3/n41 ;
   wire \add_x_22_3/n35 ;
   wire \add_x_22_3/n34 ;
   wire \add_x_22_3/n31 ;
   wire \add_x_22_3/n30 ;
   wire \add_x_22_3/n28 ;
   wire \add_x_22_3/n27 ;
   wire \add_x_22_3/n26 ;
   wire \add_x_22_3/n24 ;
   wire \add_x_22_3/n23 ;
   wire \add_x_22_3/n22 ;
   wire \add_x_22_3/n20 ;
   wire \add_x_22_3/n19 ;
   wire \add_x_22_3/n17 ;
   wire \add_x_22_3/n16 ;
   wire \add_x_22_3/n13 ;
   wire \add_x_22_3/n10 ;
   wire \add_x_22_3/n9 ;
   wire \add_x_22_3/n8 ;
   wire \add_x_22_3/n7 ;
   wire \add_x_22_3/n2 ;
   wire \add_x_22_3/n1 ;
   wire \add_x_22_2/n121 ;
   wire \add_x_22_2/n119 ;
   wire \add_x_22_2/n118 ;
   wire \add_x_22_2/n117 ;
   wire \add_x_22_2/n114 ;
   wire \add_x_22_2/n112 ;
   wire \add_x_22_2/n111 ;
   wire \add_x_22_2/n110 ;
   wire \add_x_22_2/n109 ;
   wire \add_x_22_2/n106 ;
   wire \add_x_22_2/n105 ;
   wire \add_x_22_2/n103 ;
   wire \add_x_22_2/n102 ;
   wire \add_x_22_2/n101 ;
   wire \add_x_22_2/n99 ;
   wire \add_x_22_2/n98 ;
   wire \add_x_22_2/n94 ;
   wire \add_x_22_2/n93 ;
   wire \add_x_22_2/n92 ;
   wire \add_x_22_2/n90 ;
   wire \add_x_22_2/n87 ;
   wire \add_x_22_2/n85 ;
   wire \add_x_22_2/n81 ;
   wire \add_x_22_2/n80 ;
   wire \add_x_22_2/n78 ;
   wire \add_x_22_2/n77 ;
   wire \add_x_22_2/n76 ;
   wire \add_x_22_2/n75 ;
   wire \add_x_22_2/n74 ;
   wire \add_x_22_2/n72 ;
   wire \add_x_22_2/n71 ;
   wire \add_x_22_2/n69 ;
   wire \add_x_22_2/n68 ;
   wire \add_x_22_2/n64 ;
   wire \add_x_22_2/n59 ;
   wire \add_x_22_2/n58 ;
   wire \add_x_22_2/n54 ;
   wire \add_x_22_2/n53 ;
   wire \add_x_22_2/n51 ;
   wire \add_x_22_2/n50 ;
   wire \add_x_22_2/n47 ;
   wire \add_x_22_2/n46 ;
   wire \add_x_22_2/n44 ;
   wire \add_x_22_2/n43 ;
   wire \add_x_22_2/n42 ;
   wire \add_x_22_2/n41 ;
   wire \add_x_22_2/n38 ;
   wire \add_x_22_2/n35 ;
   wire \add_x_22_2/n34 ;
   wire \add_x_22_2/n31 ;
   wire \add_x_22_2/n30 ;
   wire \add_x_22_2/n26 ;
   wire \add_x_22_2/n24 ;
   wire \add_x_22_2/n23 ;
   wire \add_x_22_2/n17 ;
   wire \add_x_22_2/n16 ;
   wire \add_x_22_2/n10 ;
   wire \add_x_22_2/n9 ;
   wire \add_x_22_2/n8 ;
   wire \add_x_22_2/n2 ;
   wire \add_x_22_2/n1 ;
   wire \add_x_22_0/n121 ;
   wire \add_x_22_0/n119 ;
   wire \add_x_22_0/n118 ;
   wire \add_x_22_0/n117 ;
   wire \add_x_22_0/n115 ;
   wire \add_x_22_0/n114 ;
   wire \add_x_22_0/n112 ;
   wire \add_x_22_0/n111 ;
   wire \add_x_22_0/n110 ;
   wire \add_x_22_0/n109 ;
   wire \add_x_22_0/n106 ;
   wire \add_x_22_0/n105 ;
   wire \add_x_22_0/n103 ;
   wire \add_x_22_0/n102 ;
   wire \add_x_22_0/n99 ;
   wire \add_x_22_0/n96 ;
   wire \add_x_22_0/n95 ;
   wire \add_x_22_0/n94 ;
   wire \add_x_22_0/n93 ;
   wire \add_x_22_0/n92 ;
   wire \add_x_22_0/n90 ;
   wire \add_x_22_0/n89 ;
   wire \add_x_22_0/n87 ;
   wire \add_x_22_0/n85 ;
   wire \add_x_22_0/n84 ;
   wire \add_x_22_0/n80 ;
   wire \add_x_22_0/n78 ;
   wire \add_x_22_0/n77 ;
   wire \add_x_22_0/n76 ;
   wire \add_x_22_0/n75 ;
   wire \add_x_22_0/n72 ;
   wire \add_x_22_0/n69 ;
   wire \add_x_22_0/n68 ;
   wire \add_x_22_0/n65 ;
   wire \add_x_22_0/n59 ;
   wire \add_x_22_0/n58 ;
   wire \add_x_22_0/n57 ;
   wire \add_x_22_0/n51 ;
   wire \add_x_22_0/n50 ;
   wire \add_x_22_0/n49 ;
   wire \add_x_22_0/n47 ;
   wire \add_x_22_0/n44 ;
   wire \add_x_22_0/n43 ;
   wire \add_x_22_0/n42 ;
   wire \add_x_22_0/n41 ;
   wire \add_x_22_0/n40 ;
   wire \add_x_22_0/n35 ;
   wire \add_x_22_0/n34 ;
   wire \add_x_22_0/n31 ;
   wire \add_x_22_0/n26 ;
   wire \add_x_22_0/n24 ;
   wire \add_x_22_0/n23 ;
   wire \add_x_22_0/n20 ;
   wire \add_x_22_0/n17 ;
   wire \add_x_22_0/n16 ;
   wire \add_x_22_0/n15 ;
   wire \add_x_22_0/n13 ;
   wire \add_x_22_0/n10 ;
   wire \add_x_22_0/n9 ;
   wire \add_x_22_0/n8 ;
   wire \add_x_22_0/n7 ;
   wire \add_x_22_0/n5 ;
   wire \add_x_22_0/n4 ;
   wire \add_x_22_0/n3 ;
   wire \add_x_22_0/n2 ;
   wire \add_x_22_0/n1 ;
   wire \DP_OP_159_297_3515/n1075 ;
   wire \DP_OP_159_297_3515/n1066 ;
   wire \DP_OP_158_296_6262/n2056 ;
   wire \DP_OP_158_296_6262/n1861 ;
   wire \DP_OP_158_296_6262/n1860 ;
   wire \add_x_19_4/n50 ;
   wire \add_x_19_4/n4 ;
   wire \add_x_19_4/n195 ;
   wire \add_x_19_4/n7 ;
   wire \add_x_19_4/n65 ;
   wire \add_x_19_4/n198 ;
   wire \add_x_19_4/n40 ;
   wire \add_x_19_4/n47 ;
   wire \add_x_19_4/n45 ;
   wire \add_x_19_4/n44 ;
   wire \add_x_19_4/n208 ;
   wire \add_x_19_4/n17 ;
   wire \add_x_19_4/n122 ;
   wire \addr_calc/fft_write_calc/counter/N48 ;
   wire \add_x_22_1/n106 ;
   wire \DP_OP_159_297_3515/n87 ;
   wire \DP_OP_159_297_3515/n85 ;
   wire \DP_OP_159_297_3515/n792 ;
   wire \DP_OP_159_297_3515/n70 ;
   wire \DP_OP_159_297_3515/n51 ;
   wire \DP_OP_159_297_3515/n5 ;
   wire \DP_OP_159_297_3515/n49 ;
   wire \DP_OP_159_297_3515/n47 ;
   wire \DP_OP_159_297_3515/n45 ;
   wire \DP_OP_159_297_3515/n3 ;
   wire \DP_OP_159_297_3515/n18 ;
   wire \DP_OP_159_297_3515/n157 ;
   wire \DP_OP_159_297_3515/n144 ;
   wire \DP_OP_159_297_3515/n142 ;
   wire \DP_OP_159_297_3515/n131 ;
   wire \DP_OP_159_297_3515/n116 ;
   wire \DP_OP_159_297_3515/n114 ;
   wire \DP_OP_159_297_3515/n112 ;
   wire \DP_OP_159_297_3515/n102 ;
   wire \DP_OP_159_297_3515/n942 ;
   wire \DP_OP_159_297_3515/n941 ;
   wire \DP_OP_159_297_3515/n861 ;
   wire \DP_OP_158_296_6262/n1891 ;
   wire \DP_OP_158_296_6262/n1883 ;
   wire \DP_OP_158_296_6262/n1882 ;
   wire \DP_OP_158_296_6262/n1906 ;
   wire \DP_OP_158_296_6262/n1878 ;
   wire \add_x_19_0/n119 ;
   wire \add_x_19_0/n117 ;
   wire \add_x_19_0/n115 ;
   wire \add_x_19_0/n114 ;
   wire \DP_OP_158_296_6262/n998 ;
   wire \DP_OP_158_296_6262/n996 ;
   wire \DP_OP_158_296_6262/n981 ;
   wire \DP_OP_158_296_6262/n962 ;
   wire \DP_OP_158_296_6262/n960 ;
   wire \DP_OP_158_296_6262/n958 ;
   wire \DP_OP_158_296_6262/n956 ;
   wire \DP_OP_158_296_6262/n948 ;
   wire \DP_OP_158_296_6262/n933 ;
   wire \DP_OP_158_296_6262/n931 ;
   wire \DP_OP_158_296_6262/n912 ;
   wire \DP_OP_158_296_6262/n899 ;
   wire \DP_OP_158_296_6262/n897 ;
   wire \DP_OP_158_296_6262/n895 ;
   wire \DP_OP_158_296_6262/n1269 ;
   wire \DP_OP_158_296_6262/n1267 ;
   wire \DP_OP_158_296_6262/n1265 ;
   wire \DP_OP_158_296_6262/n1259 ;
   wire \DP_OP_158_296_6262/n1243 ;
   wire \DP_OP_158_296_6262/n1241 ;
   wire \DP_OP_158_296_6262/n1223 ;
   wire \DP_OP_158_296_6262/n1216 ;
   wire \DP_OP_158_296_6262/n1214 ;
   wire \DP_OP_158_296_6262/n1212 ;
   wire \DP_OP_158_296_6262/n1209 ;
   wire \DP_OP_158_296_6262/n1200 ;
   wire \DP_OP_158_296_6262/n1198 ;
   wire \DP_OP_158_296_6262/n1191 ;
   wire \DP_OP_158_296_6262/n1180 ;
   wire \DP_OP_158_296_6262/n1178 ;
   wire \DP_OP_158_296_6262/n1176 ;
   wire \DP_OP_158_296_6262/n1174 ;
   wire \DP_OP_158_296_6262/n1171 ;
   wire \DP_OP_158_296_6262/n1160 ;
   wire \DP_OP_158_296_6262/n1158 ;
   wire \DP_OP_158_296_6262/n1149 ;
   wire \DP_OP_158_296_6262/n1136 ;
   wire \DP_OP_158_296_6262/n1134 ;
   wire \DP_OP_158_296_6262/n1132 ;
   wire \DP_OP_158_296_6262/n1124 ;
   wire \DP_OP_158_296_6262/n1111 ;
   wire \DP_OP_158_296_6262/n1109 ;
   wire \DP_OP_158_296_6262/n1079 ;
   wire \DP_OP_158_296_6262/n1077 ;
   wire \DP_OP_158_296_6262/n1075 ;
   wire \DP_OP_158_296_6262/n1073 ;
   wire \DP_OP_158_296_6262/n1071 ;
   wire \DP_OP_158_296_6262/n1068 ;
   wire \DP_OP_158_296_6262/n1055 ;
   wire \DP_OP_158_296_6262/n1053 ;
   wire \DP_OP_158_296_6262/n1042 ;
   wire \DP_OP_158_296_6262/n1027 ;
   wire \DP_OP_158_296_6262/n1025 ;
   wire \DP_OP_158_296_6262/n1023 ;
   wire \DP_OP_158_296_6262/n1013 ;
   wire \DP_OP_158_296_6262/n1842 ;
   wire \DP_OP_158_296_6262/n1841 ;
   wire \DP_OP_158_296_6262/n1840 ;
   wire \DP_OP_158_296_6262/n1850 ;
   wire \add_x_19_3/n9 ;
   wire \add_x_19_3/n80 ;
   wire \add_x_19_3/n200 ;
   wire \add_x_19_5/n35 ;
   wire \add_x_19_5/n34 ;
   wire \add_x_19_5/n1 ;
   wire \add_x_19_4/n161 ;
   wire \add_x_19_4/n159 ;
   wire \add_x_19_4/n158 ;
   wire \add_x_19_5/n9 ;
   wire \add_x_19_5/n80 ;
   wire \add_x_19_5/n200 ;
   wire \add_x_19_4/n80 ;
   wire \add_x_19_4/n200 ;
   wire \add_x_19_3/n138 ;
   wire \add_x_19_4/n83 ;
   wire \add_x_19_4/n92 ;
   wire \add_x_19_4/n113 ;
   wire \addr_calc/iir_write_calc/counter/N64 ;
   wire \add_x_22_5/n38 ;
   wire \addr_calc/iir_write_calc/counter/N38 ;
   wire \DP_OP_159_297_3515/n582 ;
   wire \DP_OP_159_297_3515/n569 ;
   wire \DP_OP_159_297_3515/n567 ;
   wire \DP_OP_159_297_3515/n556 ;
   wire \DP_OP_159_297_3515/n541 ;
   wire \DP_OP_159_297_3515/n539 ;
   wire \DP_OP_159_297_3515/n537 ;
   wire \DP_OP_159_297_3515/n527 ;
   wire \DP_OP_159_297_3515/n512 ;
   wire \DP_OP_159_297_3515/n510 ;
   wire \DP_OP_159_297_3515/n495 ;
   wire \DP_OP_159_297_3515/n476 ;
   wire \DP_OP_159_297_3515/n474 ;
   wire \DP_OP_159_297_3515/n472 ;
   wire \DP_OP_159_297_3515/n470 ;
   wire \DP_OP_159_297_3515/n443 ;
   wire \DP_OP_159_297_3515/n430 ;
   wire \DP_OP_159_297_3515/n428 ;
   wire \DP_OP_159_297_3515/n901 ;
   wire \DP_OP_159_297_3515/n900 ;
   wire \DP_OP_159_297_3515/n899 ;
   wire \DP_OP_159_297_3515/n903 ;
   wire \add_x_19_0/n80 ;
   wire \add_x_19_0/n200 ;
   wire \add_x_19_2/n34 ;
   wire \add_x_19_2/n1 ;
   wire \add_x_19_0/n83 ;
   wire \add_x_19_0/n92 ;
   wire \add_x_19_0/n113 ;
   wire \add_x_19_5/n99 ;
   wire \add_x_19_5/n204 ;
   wire \add_x_19_5/n13 ;
   wire \add_x_19_1/n57 ;
   wire \add_x_19_1/n5 ;
   wire \add_x_19_1/n196 ;
   wire \add_x_19_1/n71 ;
   wire \add_x_19_1/n70 ;
   wire \add_x_19_1/n180 ;
   wire \add_x_19_1/n179 ;
   wire \add_x_19_3/n180 ;
   wire \add_x_19_3/n179 ;
   wire \add_x_19_1/n170 ;
   wire \add_x_19_0/n57 ;
   wire \add_x_19_0/n196 ;
   wire \add_x_19_5/n114 ;
   wire \add_x_19_0/n77 ;
   wire \add_x_19_0/n75 ;
   wire \add_x_19_2/n47 ;
   wire \add_x_19_2/n45 ;
   wire \add_x_19_2/n44 ;
   wire \add_x_19_2/n38 ;
   wire \add_x_19_2/n43 ;
   wire \add_x_19_2/n113 ;
   wire \add_x_19_2/n136 ;
   wire \add_x_19_2/n145 ;
   wire \add_x_19_2/n157 ;
   wire \add_x_19_2/n160 ;
   wire \add_x_19_2/n162 ;
   wire \add_x_19_2/n77 ;
   wire \add_x_19_2/n75 ;
   wire \add_x_19_5/n47 ;
   wire \add_x_19_5/n45 ;
   wire \add_x_19_5/n44 ;
   wire \add_x_19_5/n77 ;
   wire \add_x_19_5/n75 ;
   wire \add_x_19_1/n9 ;
   wire \add_x_19_1/n80 ;
   wire \add_x_19_1/n200 ;
   wire \addr_calc/iir_read_calc/counter/N64 ;
   wire \add_x_22_4/n38 ;
   wire \addr_calc/iir_read_calc/counter/N38 ;
   wire \DP_OP_159_297_3515/n353 ;
   wire \DP_OP_159_297_3515/n351 ;
   wire \DP_OP_159_297_3515/n349 ;
   wire \DP_OP_159_297_3515/n343 ;
   wire \DP_OP_159_297_3515/n341 ;
   wire \DP_OP_159_297_3515/n339 ;
   wire \DP_OP_159_297_3515/n333 ;
   wire \DP_OP_159_297_3515/n317 ;
   wire \DP_OP_159_297_3515/n315 ;
   wire \DP_OP_159_297_3515/n312 ;
   wire \DP_OP_159_297_3515/n305 ;
   wire \DP_OP_159_297_3515/n303 ;
   wire \DP_OP_159_297_3515/n301 ;
   wire \DP_OP_159_297_3515/n298 ;
   wire \DP_OP_159_297_3515/n289 ;
   wire \DP_OP_159_297_3515/n287 ;
   wire \DP_OP_159_297_3515/n280 ;
   wire \DP_OP_159_297_3515/n269 ;
   wire \DP_OP_159_297_3515/n267 ;
   wire \DP_OP_159_297_3515/n265 ;
   wire \DP_OP_159_297_3515/n263 ;
   wire \DP_OP_159_297_3515/n260 ;
   wire \DP_OP_159_297_3515/n249 ;
   wire \DP_OP_159_297_3515/n247 ;
   wire \DP_OP_159_297_3515/n238 ;
   wire \DP_OP_159_297_3515/n225 ;
   wire \DP_OP_159_297_3515/n223 ;
   wire \DP_OP_159_297_3515/n221 ;
   wire \DP_OP_159_297_3515/n213 ;
   wire \DP_OP_159_297_3515/n200 ;
   wire \DP_OP_159_297_3515/n198 ;
   wire \DP_OP_159_297_3515/n185 ;
   wire \DP_OP_159_297_3515/n168 ;
   wire \DP_OP_159_297_3515/n166 ;
   wire \DP_OP_159_297_3515/n164 ;
   wire \DP_OP_159_297_3515/n162 ;
   wire \DP_OP_159_297_3515/n970 ;
   wire \DP_OP_159_297_3515/n969 ;
   wire \DP_OP_159_297_3515/n986 ;
   wire \DP_OP_159_297_3515/n985 ;
   wire \DP_OP_159_297_3515/n1041 ;
   wire \DP_OP_159_297_3515/n1040 ;
   wire \addr_calc/fir_write_calc/counter/N44 ;
   wire \add_x_22_3/n121 ;
   wire \addr_calc/fir_write_calc/counter/N50 ;
   wire \add_x_22_3/n99 ;
   wire \addr_calc/fir_write_calc/counter/N53 ;
   wire \DP_OP_158_296_6262/n1716 ;
   wire \DP_OP_158_296_6262/n1714 ;
   wire \DP_OP_158_296_6262/n1712 ;
   wire \DP_OP_158_296_6262/n1706 ;
   wire \DP_OP_158_296_6262/n1690 ;
   wire \DP_OP_158_296_6262/n1688 ;
   wire \DP_OP_158_296_6262/n1670 ;
   wire \DP_OP_158_296_6262/n1663 ;
   wire \DP_OP_158_296_6262/n1661 ;
   wire \DP_OP_158_296_6262/n1659 ;
   wire \DP_OP_158_296_6262/n1656 ;
   wire \DP_OP_158_296_6262/n1647 ;
   wire \DP_OP_158_296_6262/n1645 ;
   wire \DP_OP_158_296_6262/n1638 ;
   wire \DP_OP_158_296_6262/n1627 ;
   wire \DP_OP_158_296_6262/n1625 ;
   wire \DP_OP_158_296_6262/n1623 ;
   wire \DP_OP_158_296_6262/n1621 ;
   wire \DP_OP_158_296_6262/n1618 ;
   wire \DP_OP_158_296_6262/n1607 ;
   wire \DP_OP_158_296_6262/n1605 ;
   wire \DP_OP_158_296_6262/n1596 ;
   wire \DP_OP_158_296_6262/n1583 ;
   wire \DP_OP_158_296_6262/n1581 ;
   wire \DP_OP_158_296_6262/n1579 ;
   wire \DP_OP_158_296_6262/n1571 ;
   wire \DP_OP_158_296_6262/n1558 ;
   wire \DP_OP_158_296_6262/n1556 ;
   wire \DP_OP_158_296_6262/n1543 ;
   wire \DP_OP_158_296_6262/n1526 ;
   wire \DP_OP_158_296_6262/n1524 ;
   wire \DP_OP_158_296_6262/n1522 ;
   wire \DP_OP_158_296_6262/n1520 ;
   wire \DP_OP_158_296_6262/n1518 ;
   wire \DP_OP_158_296_6262/n1515 ;
   wire \DP_OP_158_296_6262/n1502 ;
   wire \DP_OP_158_296_6262/n1500 ;
   wire \DP_OP_158_296_6262/n1489 ;
   wire \DP_OP_158_296_6262/n1474 ;
   wire \DP_OP_158_296_6262/n1472 ;
   wire \DP_OP_158_296_6262/n1470 ;
   wire \DP_OP_158_296_6262/n1460 ;
   wire \DP_OP_158_296_6262/n1445 ;
   wire \DP_OP_158_296_6262/n1443 ;
   wire \DP_OP_158_296_6262/n1428 ;
   wire \DP_OP_158_296_6262/n1409 ;
   wire \DP_OP_158_296_6262/n1407 ;
   wire \DP_OP_158_296_6262/n1405 ;
   wire \DP_OP_158_296_6262/n1403 ;
   wire \DP_OP_158_296_6262/n1395 ;
   wire \DP_OP_158_296_6262/n1380 ;
   wire \DP_OP_158_296_6262/n1378 ;
   wire \DP_OP_158_296_6262/n1359 ;
   wire \DP_OP_158_296_6262/n1346 ;
   wire \DP_OP_158_296_6262/n1344 ;
   wire \DP_OP_158_296_6262/n1342 ;
   wire \DP_OP_158_296_6262/n1923 ;
   wire \DP_OP_158_296_6262/n1986 ;
   wire \DP_OP_158_296_6262/n1933 ;
   wire \DP_OP_158_296_6262/n1932 ;
   wire \DP_OP_158_296_6262/n1931 ;
   wire \DP_OP_158_296_6262/n1988 ;
   wire \addr_calc/fft_write_calc/counter/N61 ;
   wire \DP_OP_158_296_6262/n822 ;
   wire \DP_OP_158_296_6262/n820 ;
   wire \DP_OP_158_296_6262/n818 ;
   wire \DP_OP_158_296_6262/n812 ;
   wire \DP_OP_158_296_6262/n796 ;
   wire \DP_OP_158_296_6262/n794 ;
   wire \DP_OP_158_296_6262/n776 ;
   wire \DP_OP_158_296_6262/n769 ;
   wire \DP_OP_158_296_6262/n767 ;
   wire \DP_OP_158_296_6262/n765 ;
   wire \DP_OP_158_296_6262/n762 ;
   wire \DP_OP_158_296_6262/n753 ;
   wire \DP_OP_158_296_6262/n751 ;
   wire \DP_OP_158_296_6262/n744 ;
   wire \DP_OP_158_296_6262/n733 ;
   wire \DP_OP_158_296_6262/n731 ;
   wire \DP_OP_158_296_6262/n729 ;
   wire \DP_OP_158_296_6262/n727 ;
   wire \DP_OP_158_296_6262/n724 ;
   wire \DP_OP_158_296_6262/n713 ;
   wire \DP_OP_158_296_6262/n711 ;
   wire \DP_OP_158_296_6262/n702 ;
   wire \DP_OP_158_296_6262/n689 ;
   wire \DP_OP_158_296_6262/n687 ;
   wire \DP_OP_158_296_6262/n685 ;
   wire \DP_OP_158_296_6262/n677 ;
   wire \DP_OP_158_296_6262/n664 ;
   wire \DP_OP_158_296_6262/n662 ;
   wire \DP_OP_158_296_6262/n649 ;
   wire \DP_OP_158_296_6262/n632 ;
   wire \DP_OP_158_296_6262/n630 ;
   wire \DP_OP_158_296_6262/n628 ;
   wire \DP_OP_158_296_6262/n626 ;
   wire \DP_OP_158_296_6262/n621 ;
   wire \DP_OP_158_296_6262/n608 ;
   wire \DP_OP_158_296_6262/n606 ;
   wire \DP_OP_158_296_6262/n595 ;
   wire \DP_OP_158_296_6262/n580 ;
   wire \DP_OP_158_296_6262/n578 ;
   wire \DP_OP_158_296_6262/n576 ;
   wire \DP_OP_158_296_6262/n566 ;
   wire \DP_OP_158_296_6262/n549 ;
   wire \DP_OP_158_296_6262/n534 ;
   wire \DP_OP_158_296_6262/n515 ;
   wire \DP_OP_158_296_6262/n513 ;
   wire \DP_OP_158_296_6262/n511 ;
   wire \DP_OP_158_296_6262/n509 ;
   wire \DP_OP_158_296_6262/n501 ;
   wire \DP_OP_158_296_6262/n486 ;
   wire \DP_OP_158_296_6262/n484 ;
   wire \DP_OP_158_296_6262/n465 ;
   wire \DP_OP_158_296_6262/n452 ;
   wire \DP_OP_158_296_6262/n450 ;
   wire \DP_OP_158_296_6262/n1889 ;
   wire \DP_OP_158_296_6262/n1888 ;
   wire \DP_OP_159_297_3515/n1014 ;
   wire \addr_calc/iir_read_calc/counter/N47 ;
   wire \addr_calc/iir_read_calc/counter/N49 ;
   wire \addr_calc/fir_write_calc/counter/N58 ;
   wire \add_x_22_3/n65 ;
   wire \add_x_19_2/n50 ;
   wire \add_x_19_2/n4 ;
   wire \add_x_19_2/n195 ;
   wire \add_x_19_2/n7 ;
   wire \add_x_19_2/n65 ;
   wire \add_x_19_2/n198 ;
   wire \add_x_19_2/n71 ;
   wire \add_x_19_2/n70 ;
   wire \add_x_19_2/n119 ;
   wire \add_x_19_2/n117 ;
   wire \add_x_19_2/n115 ;
   wire \add_x_19_2/n114 ;
   wire \addr_calc/fir_read_calc/counter/N58 ;
   wire \add_x_22_2/n65 ;
   wire \addr_calc/iir_write_calc/counter/N63 ;
   wire \add_x_19_1/n99 ;
   wire \add_x_19_1/n204 ;
   wire \add_x_19_1/n13 ;
   wire \addr_calc/fft_write_calc/counter/N69 ;
   wire \add_x_19_1/n119 ;
   wire \add_x_19_1/n117 ;
   wire \add_x_19_1/n115 ;
   wire \add_x_19_1/n114 ;
   wire \add_x_19_1/n161 ;
   wire \add_x_19_1/n159 ;
   wire \add_x_19_1/n158 ;
   wire \add_x_19_1/n83 ;
   wire \add_x_19_1/n157 ;
   wire \add_x_19_1/n169 ;
   wire \add_x_19_1/n92 ;
   wire \add_x_19_1/n113 ;
   wire \add_x_19_1/n171 ;
   wire n1137;
   wire n1138;
   wire n1140;
   wire n1141;
   wire n1142;
   wire n1143;
   wire n1146;
   wire n1147;
   wire n1149;
   wire n1150;
   wire n1153;
   wire n1154;
   wire n1155;
   wire n1156;
   wire n1157;
   wire n1158;
   wire n1159;
   wire n1160;
   wire n1161;
   wire n1162;
   wire n1163;
   wire n1164;
   wire n1166;
   wire n1167;
   wire n1168;
   wire n1169;
   wire n1170;
   wire n1171;
   wire n1172;
   wire n1174;
   wire n1175;
   wire n1176;
   wire n1177;
   wire n1178;
   wire n1179;
   wire n1180;
   wire n1181;
   wire n1182;
   wire n1184;
   wire n1185;
   wire n1186;
   wire n1187;
   wire n1188;
   wire n1189;
   wire n1190;
   wire n1191;
   wire n1192;
   wire n1194;
   wire n1195;
   wire n1196;
   wire n1197;
   wire n1198;
   wire n1199;
   wire n1200;
   wire n1201;
   wire n1202;
   wire n1203;
   wire n1204;
   wire n1206;
   wire n1207;
   wire n1208;
   wire n1209;
   wire n1210;
   wire n1211;
   wire n1212;
   wire n1213;
   wire n1214;
   wire n1215;
   wire n1216;
   wire n1217;
   wire n1218;
   wire n1220;
   wire n1221;
   wire n1223;
   wire n1224;
   wire n1225;
   wire n1226;
   wire n1227;
   wire n1228;
   wire n1229;
   wire n1230;
   wire n1231;
   wire n1232;
   wire n1233;
   wire n1234;
   wire n1235;
   wire n1236;
   wire n1237;
   wire n1238;
   wire n1239;
   wire n1240;
   wire n1241;
   wire n1242;
   wire n1243;
   wire n1245;
   wire n1246;
   wire n1247;
   wire n1248;
   wire n1249;
   wire n1250;
   wire n1251;
   wire n1252;
   wire n1253;
   wire n1254;
   wire n1255;
   wire n1272;
   wire n1273;
   wire n1274;
   wire n1275;
   wire n1276;
   wire n1277;
   wire n1278;
   wire n1279;
   wire n1280;
   wire n1281;
   wire n1282;
   wire n1283;
   wire n1284;
   wire n1285;
   wire n1286;
   wire n1287;
   wire n1288;
   wire n1289;
   wire n1290;
   wire n1291;
   wire n1292;
   wire n1293;
   wire n1294;
   wire n1295;
   wire n1296;
   wire n1297;
   wire n1298;
   wire n1299;
   wire n1300;
   wire n1301;
   wire n1302;
   wire n1303;
   wire n1304;
   wire n1305;
   wire n1306;
   wire n1307;
   wire n1308;
   wire n1309;
   wire n1310;
   wire n1311;
   wire n1312;
   wire n1314;
   wire n1315;
   wire n1316;
   wire n1317;
   wire n1318;
   wire n1319;
   wire n1321;
   wire n1322;
   wire n1323;
   wire n1324;
   wire n1325;
   wire n1326;
   wire n1327;
   wire n1328;
   wire n1329;
   wire n1330;
   wire n1331;
   wire n1332;
   wire n1333;
   wire n1334;
   wire n1335;
   wire n1336;
   wire n1337;
   wire n1338;
   wire n1339;
   wire n1340;
   wire n1341;
   wire n1342;
   wire n1343;
   wire n1344;
   wire n1345;
   wire n1346;
   wire n1347;
   wire n1348;
   wire n1349;
   wire n1350;
   wire n1351;
   wire n1352;
   wire n1353;
   wire n1354;
   wire n1355;
   wire n1356;
   wire n1357;
   wire n1358;
   wire n1359;
   wire n1360;
   wire n1361;
   wire n1362;
   wire n1363;
   wire n1364;
   wire n1365;
   wire n1366;
   wire n1367;
   wire n1368;
   wire n1369;
   wire n1370;
   wire n1371;
   wire n1372;
   wire n1373;
   wire n1374;
   wire n1375;
   wire n1376;
   wire n1377;
   wire n1378;
   wire n1379;
   wire n1380;
   wire n1381;
   wire n1382;
   wire n1383;
   wire n1384;
   wire n1385;
   wire n1386;
   wire n1387;
   wire n1388;
   wire n1389;
   wire n1390;
   wire n1391;
   wire n1392;
   wire n1393;
   wire n1394;
   wire n1395;
   wire n1396;
   wire n1397;
   wire n1398;
   wire n1399;
   wire n1400;
   wire n1401;
   wire n1402;
   wire n1403;
   wire n1404;
   wire n1405;
   wire n1406;
   wire n1407;
   wire n1408;
   wire n1409;
   wire n1410;
   wire n1412;
   wire n1414;
   wire n1415;
   wire n1416;
   wire n1417;
   wire n1418;
   wire n1419;
   wire n1420;
   wire n1421;
   wire n1422;
   wire n1423;
   wire n1424;
   wire n1425;
   wire n1426;
   wire n1427;
   wire n1428;
   wire n1429;
   wire n1430;
   wire n1431;
   wire n1432;
   wire n1433;
   wire n1434;
   wire n1435;
   wire n1436;
   wire n1437;
   wire n1438;
   wire n1439;
   wire n1440;
   wire n1441;
   wire n1442;
   wire n1443;
   wire n1444;
   wire n1445;
   wire n1446;
   wire n1447;
   wire n1448;
   wire n1449;
   wire n1450;
   wire n1451;
   wire n1452;
   wire n1453;
   wire n1454;
   wire n1455;
   wire n1459;
   wire n1461;
   wire n1462;
   wire n1463;
   wire n1464;
   wire n1465;
   wire n1466;
   wire n1467;
   wire n1468;
   wire n1469;
   wire n1470;
   wire n1471;
   wire n1478;
   wire n1479;
   wire n1532;
   wire n1533;
   wire n1534;
   wire n1536;
   wire n1537;
   wire n1538;
   wire n1539;
   wire n1540;
   wire n1541;
   wire n1542;
   wire n1543;
   wire n1544;
   wire n1545;
   wire n1546;
   wire n1547;
   wire n1548;
   wire n1549;
   wire n1550;
   wire n1551;
   wire n1552;
   wire n1553;
   wire n1554;
   wire n1555;
   wire n1556;
   wire n1557;
   wire n1558;
   wire n1560;
   wire n1561;
   wire n1563;
   wire n1564;
   wire n1565;
   wire n1566;
   wire n1567;
   wire n1568;
   wire n1569;
   wire n1570;
   wire n1571;
   wire n1572;
   wire n1573;
   wire n1574;
   wire n1575;
   wire n1576;
   wire n1577;
   wire n1578;
   wire n1583;
   wire n1584;
   wire n1585;
   wire n1586;
   wire n1587;
   wire n1588;
   wire n1589;
   wire n1590;
   wire n1591;
   wire n1592;
   wire n1593;
   wire n1594;
   wire n1595;
   wire n1596;
   wire n1597;
   wire n1598;
   wire n1599;
   wire n1600;
   wire n1601;
   wire n1602;
   wire n1603;
   wire n1604;
   wire n1605;
   wire n1606;
   wire n1607;
   wire n1608;
   wire n1609;
   wire n1611;
   wire n1612;
   wire n1613;
   wire n1615;
   wire n1616;
   wire n1617;
   wire n1618;
   wire n1619;
   wire n1620;
   wire n1621;
   wire n1622;
   wire n1623;
   wire n1624;
   wire n1625;
   wire n1626;
   wire n1627;
   wire n1628;
   wire n1629;
   wire n1630;
   wire n1631;
   wire n1632;
   wire n1633;
   wire n1634;
   wire n1635;
   wire n1636;
   wire n1637;
   wire n1638;
   wire n1639;
   wire n1640;
   wire n1641;
   wire n1642;
   wire n1643;
   wire n1644;
   wire n1645;
   wire n1646;
   wire n1647;
   wire n1651;
   wire n1652;
   wire n1653;
   wire n1654;
   wire n1655;
   wire n1656;
   wire n1657;
   wire n1658;
   wire n1659;
   wire n1660;
   wire n1661;
   wire n1662;
   wire n1664;
   wire n1665;
   wire n1666;
   wire n1667;
   wire n1668;
   wire n1670;
   wire n1675;
   wire n1677;
   wire n1678;
   wire n1679;
   wire n1680;
   wire n1681;
   wire n1682;
   wire n1683;
   wire n1685;
   wire n1686;
   wire n1687;
   wire n1688;
   wire n1689;
   wire n1690;
   wire n1691;
   wire n1692;
   wire n1693;
   wire n1696;
   wire n1697;
   wire n1698;
   wire n1699;
   wire n1701;
   wire n1702;
   wire n1703;
   wire n1715;
   wire n1716;
   wire n1717;
   wire n1718;
   wire n1728;
   wire n1729;
   wire n1730;
   wire n1731;
   wire n1732;
   wire n1733;
   wire n1734;
   wire n1735;
   wire n1736;
   wire n1737;
   wire n1738;
   wire n1740;
   wire n1751;
   wire n1754;
   wire n1755;
   wire n1756;
   wire n1758;
   wire n1762;
   wire n1763;
   wire n1775;
   wire n1776;
   wire n1778;
   wire n1779;
   wire n1780;
   wire n1781;
   wire n1782;
   wire n1784;
   wire n1785;
   wire n1787;
   wire n1788;
   wire n1789;
   wire n1792;
   wire n1797;
   wire n1818;
   wire n1828;
   wire n1829;
   wire n1830;
   wire n1834;
   wire n1835;
   wire n1837;
   wire n1838;
   wire n1839;
   wire n1840;
   wire n1841;
   wire n1842;
   wire n1850;
   wire n1851;
   wire n1852;
   wire n1853;
   wire n1860;
   wire n1861;
   wire n1866;
   wire n1867;
   wire n1869;
   wire n1870;
   wire n1871;
   wire n1872;
   wire n1874;
   wire n1875;
   wire n1876;
   wire n1877;
   wire n1878;
   wire n1879;
   wire n1880;
   wire n1881;
   wire n1882;
   wire n1883;
   wire n1884;
   wire n1885;
   wire n1886;
   wire n1887;
   wire n1888;
   wire n1889;
   wire n1890;
   wire n1891;
   wire n1892;
   wire n1893;
   wire n1895;
   wire n1896;
   wire n1897;
   wire n1898;
   wire n1899;
   wire n1900;
   wire n1901;
   wire n1902;
   wire n1906;
   wire n1907;
   wire n1908;
   wire n1912;
   wire n1913;
   wire n1914;
   wire n1915;
   wire n1916;
   wire n1917;
   wire n1918;
   wire n1919;
   wire n1920;
   wire n1921;
   wire n1922;
   wire n1923;
   wire n1924;
   wire n1925;
   wire n1926;
   wire n1927;
   wire n1930;
   wire n1931;
   wire n1932;
   wire n1934;
   wire n1935;
   wire n1936;
   wire n1937;
   wire n1938;
   wire n1939;
   wire n1940;
   wire n1941;
   wire n1942;
   wire n1943;
   wire n1944;
   wire n1945;
   wire n1946;
   wire n1947;
   wire n1949;
   wire n1950;
   wire n1951;
   wire n1954;
   wire n1955;
   wire n1956;
   wire n1957;
   wire n1958;
   wire n1961;
   wire n1962;
   wire n1963;
   wire n1964;
   wire n1965;
   wire n1966;
   wire n1967;
   wire n1968;
   wire n1969;
   wire n1970;
   wire n1971;
   wire n1972;
   wire n1973;
   wire n1974;
   wire n1975;
   wire n1976;
   wire n1978;
   wire n1979;
   wire n1981;
   wire n1982;
   wire n1983;
   wire n1984;
   wire n1985;
   wire n1987;
   wire n1988;
   wire n1989;
   wire n1990;
   wire n1991;
   wire n1994;
   wire n1997;
   wire n2001;
   wire n2002;
   wire n2003;
   wire n2004;
   wire n2005;
   wire n2006;
   wire n2007;
   wire n2012;
   wire n2015;
   wire n2018;
   wire n2019;
   wire n2020;
   wire n2023;
   wire n2024;
   wire n2025;
   wire n2026;
   wire n2027;
   wire n2028;
   wire n2031;
   wire n2032;
   wire n2033;
   wire n2034;
   wire n2036;
   wire n2037;
   wire n2038;
   wire n2039;
   wire n2040;
   wire n2041;
   wire n2042;
   wire n2043;
   wire n2044;
   wire n2045;
   wire n2046;
   wire n2047;
   wire n2048;
   wire n2049;
   wire n2050;
   wire n2051;
   wire n2056;
   wire n2057;
   wire n2058;
   wire n2060;
   wire n2061;
   wire n2062;
   wire n2063;
   wire n2065;
   wire n2066;
   wire n2070;
   wire n2071;
   wire n2072;
   wire n2073;
   wire n2074;
   wire n2093;
   wire n2108;
   wire n2311;
   wire n2324;
   wire n2325;
   wire n2330;
   wire n2341;
   wire n2343;
   wire n2345;
   wire n2346;
   wire n2347;
   wire n2348;
   wire n2349;
   wire n2350;
   wire n2351;
   wire n2352;
   wire n2353;
   wire n2354;
   wire n2355;
   wire n2356;
   wire n2357;
   wire n2358;
   wire n2359;
   wire n2360;
   wire n2362;
   wire n2364;
   wire n2365;
   wire n2366;
   wire n2367;
   wire n2368;
   wire n2369;
   wire n2371;
   wire n2372;
   wire n2441;
   wire n2501;
   wire n2502;
   wire n2503;
   wire n2504;
   wire n2505;
   wire n2506;
   wire n2507;
   wire n2508;
   wire n2509;
   wire n2510;
   wire n2511;
   wire n2512;
   wire n2513;
   wire n2514;
   wire n2515;
   wire n2516;
   wire n2517;
   wire n2518;
   wire n2519;
   wire n2520;
   wire n2521;
   wire n2522;
   wire n2523;
   wire n2524;
   wire n2525;
   wire n2526;
   wire n2527;
   wire n2528;
   wire n2529;
   wire n2530;
   wire n2531;
   wire n2532;
   wire n2533;
   wire n2534;
   wire n2535;
   wire n2536;
   wire n2537;
   wire n2538;
   wire n2539;
   wire n2540;
   wire n2541;
   wire n2542;
   wire n2543;
   wire n2544;
   wire n2545;
   wire n2546;
   wire n2547;
   wire n2548;
   wire n2553;
   wire n2554;
   wire n2555;
   wire n2556;
   wire n2557;
   wire n2558;
   wire n2559;
   wire n2560;
   wire n2561;
   wire n2562;
   wire n2563;
   wire n2564;
   wire n2565;
   wire n2566;
   wire n2567;
   wire n2568;
   wire n2569;
   wire n2570;
   wire n2572;
   wire n2573;
   wire n2574;
   wire n2575;
   wire n2577;
   wire n2578;
   wire n2579;
   wire n2580;
   wire n2583;
   wire n2585;
   wire n2587;
   wire n2588;
   wire n2589;
   wire n2590;
   wire n2591;
   wire n2592;
   wire n2593;
   wire n2594;
   wire n2595;
   wire n2596;
   wire n2597;
   wire n2598;
   wire n2599;
   wire n2600;
   wire n2601;
   wire n2602;
   wire n2603;
   wire n2604;
   wire n2605;
   wire n2606;
   wire n2607;
   wire n2608;
   wire n2609;
   wire n2610;
   wire n2611;
   wire n2612;
   wire n2613;
   wire n2614;
   wire n2615;
   wire n2616;
   wire n2617;
   wire n2618;
   wire n2619;
   wire n2620;
   wire n2621;
   wire n2622;
   wire n2623;
   wire n2624;
   wire n2625;
   wire n2626;
   wire n2627;
   wire n2628;
   wire n2629;
   wire n2630;
   wire n2631;
   wire n2632;
   wire n2633;
   wire n2634;
   wire n2641;
   wire n2642;
   wire n2643;
   wire n2644;
   wire n2645;
   wire n2646;
   wire n2654;
   wire n2783;
   wire n2784;
   wire n2785;
   wire n2786;
   wire n2787;
   wire n2788;
   wire n2789;
   wire n2790;
   wire n2791;
   wire n2792;
   wire n2793;
   wire n2794;
   wire n2795;
   wire n2796;
   wire n2797;
   wire n2798;
   wire n2799;
   wire n2800;
   wire n2801;
   wire n2802;
   wire n2803;
   wire n2804;
   wire n2805;
   wire n2806;
   wire n2807;
   wire n2808;
   wire n2809;
   wire n2810;
   wire n2811;
   wire n2812;
   wire n2813;

   CLKINVX16TS clk__L1_I0 (.Y(clk__L1_N0), 
	.A(clk));
   BUFX3TS FE_OCP_RBC1982_add_x_19_4_n157 (.Y(FE_OCP_RBN1982_add_x_19_4_n157), 
	.A(FE_OCP_RBN1981_add_x_19_4_n157));
   BUFX16TS FE_OCP_RBC1981_add_x_19_4_n157 (.Y(FE_OCP_RBN1981_add_x_19_4_n157), 
	.A(\add_x_19_4/n157 ));
   BUFX4TS FE_OCP_RBC1980_add_x_19_4_n178 (.Y(FE_OCP_RBN1980_add_x_19_4_n178), 
	.A(\add_x_19_4/n178 ));
   BUFX3TS FE_OCP_RBC1979_add_x_19_4_n178 (.Y(FE_OCP_RBN1979_add_x_19_4_n178), 
	.A(FE_OCP_RBN1980_add_x_19_4_n178));
   INVX3TS FE_OCP_RBC1978_add_x_19_4_n178 (.Y(FE_OCP_RBN1978_add_x_19_4_n178), 
	.A(FE_OCP_RBN1980_add_x_19_4_n178));
   BUFX20TS FE_OCP_RBC1974_offset_1_ (.Y(FE_OCP_RBN1974_offset_1_), 
	.A(offset[1]));
   BUFX20TS FE_OCP_RBC1973_offset_1_ (.Y(FE_OCP_RBN1973_offset_1_), 
	.A(FE_OCP_RBN1974_offset_1_));
   BUFX20TS FE_OCP_DRV_C1968_filesize_8_ (.Y(FE_OCP_DRV_N1968_filesize_8_), 
	.A(filesize[8]));
   INVX2TS FE_RC_1088_0 (.Y(FE_RN_468_0), 
	.A(\add_x_19_4/n72 ));
   INVX4TS FE_RC_1087_0 (.Y(FE_RN_467_0), 
	.A(\add_x_19_4/n73 ));
   OAI21X4TS FE_RC_1086_0 (.Y(\add_x_19_4/n69 ), 
	.B0(FE_RN_467_0), 
	.A1(FE_RN_468_0), 
	.A0(FE_OFN527_add_x_19_4_n113));
   NOR2X2TS FE_RC_1076_0 (.Y(FE_RN_459_0), 
	.B(\add_x_19_4/n184 ), 
	.A(\add_x_19_4/n181 ));
   OAI21X2TS FE_RC_1075_0 (.Y(FE_RN_458_0), 
	.B0(\add_x_19_4/n182 ), 
	.A1(\add_x_19_4/n185 ), 
	.A0(\add_x_19_4/n181 ));
   AOI21X4TS FE_RC_1074_0 (.Y(\add_x_19_4/n178 ), 
	.B0(FE_RN_458_0), 
	.A1(FE_RN_459_0), 
	.A0(\add_x_19_4/n187 ));
   AOI21X4TS FE_RC_1072_0 (.Y(\add_x_19_5/n94 ), 
	.B0(\add_x_19_5/n96 ), 
	.A1(\add_x_19_5/n95 ), 
	.A0(\add_x_19_5/n104 ));
   OAI21X2TS FE_RC_1071_0 (.Y(\add_x_19_3/n180 ), 
	.B0(\add_x_19_3/n182 ), 
	.A1(\add_x_19_3/n181 ), 
	.A0(\add_x_19_3/n185 ));
   CLKINVX2TS FE_RC_1052_0 (.Y(\add_x_19_2/n178 ), 
	.A(FE_RN_444_0));
   INVX2TS FE_RC_1051_0 (.Y(FE_RN_450_0), 
	.A(FE_RN_173_0));
   NOR2X4TS FE_RC_1050_0 (.Y(FE_RN_449_0), 
	.B(FE_RN_175_0), 
	.A(FE_RN_174_0));
   NOR2X2TS FE_RC_1049_0 (.Y(FE_RN_448_0), 
	.B(FE_RN_450_0), 
	.A(FE_RN_449_0));
   INVX2TS FE_RC_1048_0 (.Y(FE_RN_447_0), 
	.A(FE_RN_176_0));
   INVX2TS FE_RC_1047_0 (.Y(FE_RN_446_0), 
	.A(n1548));
   NAND2X2TS FE_RC_1046_0 (.Y(FE_RN_445_0), 
	.B(n1547), 
	.A(\add_x_19_2/n187 ));
   NAND2X2TS FE_RC_1045_0 (.Y(FE_RN_444_0), 
	.B(FE_RN_446_0), 
	.A(FE_RN_445_0));
   NAND2X2TS FE_RC_1044_0 (.Y(FE_RN_443_0), 
	.B(FE_RN_447_0), 
	.A(FE_RN_444_0));
   NAND2X2TS FE_RC_1043_0 (.Y(\add_x_19_2/n157 ), 
	.B(FE_RN_448_0), 
	.A(FE_RN_443_0));
   BUFX20TS FE_RC_1036_0 (.Y(FE_OFN402_offset_14_), 
	.A(offset[14]));
   BUFX20TS FE_RC_1035_0 (.Y(FE_OFN404_offset_14_), 
	.A(offset[14]));
   INVX2TS FE_RC_1034_0 (.Y(FE_RN_438_0), 
	.A(n2003));
   NAND2BX4TS FE_RC_1033_0 (.Y(n1545), 
	.B(FE_RN_438_0), 
	.AN(offset[14]));
   BUFX20TS FE_RC_1032_0 (.Y(FE_OCPUNCON1873_offset_11_), 
	.A(offset[11]));
   BUFX20TS FE_RC_1031_0 (.Y(FE_OCPN1905_FE_OCPUNCON1873_offset_11_), 
	.A(offset[11]));
   BUFX20TS FE_RC_1030_0 (.Y(FE_OFN390_offset_17_), 
	.A(offset[17]));
   BUFX20TS FE_RC_1028_0 (.Y(FE_OFN426_offset_8_), 
	.A(offset[8]));
   NAND2X1TS FE_RC_1021_0 (.Y(\add_x_19_3/n93 ), 
	.B(\add_x_19_3/n95 ), 
	.A(\add_x_19_3/n103 ));
   NAND2X2TS FE_RC_1020_0 (.Y(FE_RN_437_0), 
	.B(\add_x_19_3/n95 ), 
	.A(\add_x_19_3/n103 ));
   NOR2X2TS FE_RC_1019_0 (.Y(\add_x_19_3/n72 ), 
	.B(\add_x_19_3/n74 ), 
	.A(FE_RN_437_0));
   BUFX3TS FE_OCP_RBC1957_FE_OFN520_add_x_19_1_n157 (.Y(FE_OCP_RBN1957_FE_OFN520_add_x_19_1_n157), 
	.A(FE_OCP_RBN1956_FE_OFN520_add_x_19_1_n157));
   INVX6TS FE_OCP_RBC1956_FE_OFN520_add_x_19_1_n157 (.Y(FE_OCP_RBN1956_FE_OFN520_add_x_19_1_n157), 
	.A(FE_OFN520_add_x_19_1_n157));
   INVX1TS FE_OCP_RBC1955_add_x_19_1_n187 (.Y(FE_OCP_RBN1955_add_x_19_1_n187), 
	.A(\add_x_19_1/n187 ));
   BUFX12TS FE_OCPC1947_n1149 (.Y(FE_OCPN1947_n1149), 
	.A(n1149));
   BUFX8TS FE_OCPC1945_offset_2_ (.Y(FE_OCPN1945_offset_2_), 
	.A(FE_OCPN1944_offset_2_));
   BUFX8TS FE_OCPC1944_offset_2_ (.Y(FE_OCPN1944_offset_2_), 
	.A(offset[2]));
   NAND2X4TS FE_RC_1012_0 (.Y(FE_RN_431_0), 
	.B(n1584), 
	.A(FE_OCPUNCON1650_add_x_19_4_n43));
   NAND2X4TS FE_RC_1011_0 (.Y(n1356), 
	.B(n1585), 
	.A(FE_RN_431_0));
   AOI21X4TS FE_RC_1007_0 (.Y(\add_x_19_1/n136 ), 
	.B0(n1272), 
	.A1(\add_x_19_1/n150 ), 
	.A0(\add_x_19_1/n137 ));
   OAI22X4TS FE_RC_990_0 (.Y(\add_x_19_2/n38 ), 
	.B1(n2633), 
	.B0(FE_RN_157_0), 
	.A1(FE_RN_157_0), 
	.A0(\add_x_19_2/n43 ));
   INVX2TS FE_RC_989_0 (.Y(FE_RN_420_0), 
	.A(\add_x_19_2/n36 ));
   NAND2X2TS FE_RC_988_0 (.Y(FE_RN_419_0), 
	.B(FE_RN_420_0), 
	.A(FE_RN_157_0));
   NAND2X2TS FE_RC_987_0 (.Y(FE_RN_418_0), 
	.B(\add_x_19_2/n37 ), 
	.A(FE_RN_419_0));
   NAND2X2TS FE_RC_986_0 (.Y(FE_RN_417_0), 
	.B(\add_x_19_2/n1 ), 
	.A(FE_RN_418_0));
   INVX2TS FE_RC_985_0 (.Y(FE_RN_416_0), 
	.A(\add_x_19_2/n1 ));
   INVX2TS FE_RC_984_0 (.Y(FE_RN_415_0), 
	.A(\add_x_19_2/n36 ));
   OAI21X2TS FE_RC_983_0 (.Y(FE_RN_414_0), 
	.B0(FE_RN_415_0), 
	.A1(FE_RN_157_0), 
	.A0(n2633));
   NAND3X2TS FE_RC_982_0 (.Y(FE_RN_413_0), 
	.C(FE_RN_416_0), 
	.B(\add_x_19_2/n37 ), 
	.A(FE_RN_414_0));
   INVX2TS FE_RC_981_0 (.Y(FE_RN_412_0), 
	.A(\add_x_19_2/n36 ));
   NAND4X4TS FE_RC_980_0 (.Y(FE_RN_411_0), 
	.D(\add_x_19_2/n1 ), 
	.C(FE_RN_412_0), 
	.B(n2633), 
	.A(\add_x_19_2/n43 ));
   INVX2TS FE_RC_979_0 (.Y(FE_RN_410_0), 
	.A(FE_RN_157_0));
   NAND4BBX4TS FE_RC_978_0 (.Y(FE_RN_409_0), 
	.D(FE_RN_410_0), 
	.C(\add_x_19_2/n37 ), 
	.BN(\add_x_19_2/n1 ), 
	.AN(\add_x_19_2/n43 ));
   NAND4X4TS FE_RC_977_0 (.Y(\addr_calc/fir_read_addr[31] ), 
	.D(FE_RN_417_0), 
	.C(FE_RN_413_0), 
	.B(FE_RN_411_0), 
	.A(FE_RN_409_0));
   BUFX12TS FE_RC_974_0 (.Y(FE_OCPUNCON1565_n1789), 
	.A(n1789));
   BUFX8TS FE_RC_973_0 (.Y(FE_OCPUNCON1566_n1789), 
	.A(n1789));
   BUFX6TS FE_RC_952_0 (.Y(FE_OFN112_DP_OP_158_296_6262_n1791), 
	.A(\DP_OP_158_296_6262/n1791 ));
   BUFX6TS FE_RC_951_0 (.Y(FE_OFN113_DP_OP_158_296_6262_n1791), 
	.A(\DP_OP_158_296_6262/n1791 ));
   BUFX20TS FE_RC_912_0 (.Y(FE_OFN403_offset_14_), 
	.A(offset[14]));
   BUFX20TS FE_RC_911_0 (.Y(FE_OFN405_offset_14_), 
	.A(offset[14]));
   NOR2X8TS FE_RC_910_0 (.Y(\add_x_19_5/n123 ), 
	.B(\addr_calc/iir_write_calc/count[14] ), 
	.A(offset[14]));
   BUFX20TS FE_RC_909_0 (.Y(FE_OCPUNCON1563_offset_3_), 
	.A(offset[3]));
   BUFX20TS FE_RC_908_0 (.Y(FE_OFN449_offset_3_), 
	.A(offset[3]));
   NOR2X8TS FE_RC_907_0 (.Y(\add_x_19_3/n181 ), 
	.B(\addr_calc/fir_write_calc/count[3] ), 
	.A(offset[3]));
   BUFX20TS FE_RC_906_0 (.Y(FE_OCPUNCON1684_offset_6_), 
	.A(offset[6]));
   BUFX20TS FE_RC_905_0 (.Y(FE_OFN436_offset_6_), 
	.A(offset[6]));
   NAND2X8TS FE_RC_904_0 (.Y(\add_x_19_5/n166 ), 
	.B(offset[6]), 
	.A(\addr_calc/iir_write_calc/count[6] ));
   BUFX20TS FE_RC_903_0 (.Y(FE_OCPUNCON1066_offset_3_), 
	.A(offset[3]));
   BUFX20TS FE_RC_902_0 (.Y(FE_OCPN1904_FE_OCPUNCON1066_offset_3_), 
	.A(offset[3]));
   BUFX20TS FE_RC_901_0 (.Y(FE_OCPUNCON1940_offset_15_), 
	.A(offset[15]));
   BUFX20TS FE_RC_900_0 (.Y(FE_OFN399_offset_15_), 
	.A(offset[15]));
   BUFX20TS FE_OCPUNCOC1943_FE_OFN407_offset_13_ (.Y(FE_OCPUNCON1943_FE_OFN407_offset_13_), 
	.A(FE_OFN407_offset_13_));
   BUFX12TS FE_OCPUNCOC1942_FE_OFN399_offset_15_ (.Y(FE_OCPUNCON1942_FE_OFN399_offset_15_), 
	.A(FE_OFN399_offset_15_));
   BUFX20TS FE_OCPUNCOC1941_offset_13_ (.Y(FE_OCPUNCON1941_offset_13_), 
	.A(offset[13]));
   NAND2X2TS FE_RC_897_0 (.Y(FE_RN_371_0), 
	.B(n1867), 
	.A(FE_OCPUNCON1093_n2805));
   OAI2BB1X2TS FE_RC_896_0 (.Y(n1125), 
	.B0(FE_RN_371_0), 
	.A1N(FE_OFN51_n2803), 
	.A0N(\addr_calc/fir_write_calc/counter/N48 ));
   OAI21X4TS FE_RC_891_0 (.Y(\add_x_19_4/n73 ), 
	.B0(\add_x_19_4/n75 ), 
	.A1(\add_x_19_4/n74 ), 
	.A0(\add_x_19_4/n94 ));
   AOI21X2TS FE_RC_889_0 (.Y(\add_x_19_2/n94 ), 
	.B0(\add_x_19_2/n96 ), 
	.A1(\add_x_19_2/n104 ), 
	.A0(\add_x_19_2/n95 ));
   AOI21X4TS FE_RC_888_0 (.Y(\add_x_19_0/n136 ), 
	.B0(FE_RN_99_0), 
	.A1(\add_x_19_0/n150 ), 
	.A0(\add_x_19_0/n137 ));
   AOI21X4TS FE_RC_887_0 (.Y(\add_x_19_3/n178 ), 
	.B0(\add_x_19_3/n180 ), 
	.A1(\add_x_19_3/n187 ), 
	.A0(\add_x_19_3/n179 ));
   OAI21X2TS FE_RC_886_0 (.Y(FE_RN_105_0), 
	.B0(\add_x_19_5/n163 ), 
	.A1(\add_x_19_5/n162 ), 
	.A0(\add_x_19_5/n166 ));
   OAI21X2TS FE_RC_885_0 (.Y(\add_x_19_5/n138 ), 
	.B0(\add_x_19_5/n140 ), 
	.A1(\add_x_19_5/n145 ), 
	.A0(\add_x_19_5/n139 ));
   OAI21X2TS FE_RC_882_0 (.Y(n1272), 
	.B0(\add_x_19_1/n140 ), 
	.A1(\add_x_19_1/n145 ), 
	.A0(\add_x_19_1/n139 ));
   OAI21X2TS FE_RC_881_0 (.Y(\add_x_19_2/n187 ), 
	.B0(\add_x_19_2/n189 ), 
	.A1(\add_x_19_2/n191 ), 
	.A0(\add_x_19_2/n188 ));
   INVX12TS FE_OCP_RBC1925_add_x_19_4_n157 (.Y(FE_OCP_RBN1925_add_x_19_4_n157), 
	.A(FE_OCP_RBN1982_add_x_19_4_n157));
   BUFX20TS FE_OCP_RBC1919_offset_1_ (.Y(FE_OCP_RBN1919_offset_1_), 
	.A(FE_OCP_RBN1973_offset_1_));
   CLKBUFX2TS FE_OCPC1911_FE_OFN17_n2797 (.Y(FE_OCPN1911_FE_OFN17_n2797), 
	.A(FE_OFN17_n2797));
   BUFX2TS FE_OCPC1910_n1736 (.Y(FE_OCPN1910_n1736), 
	.A(n1736));
   CLKBUFX2TS FE_OCPC1908_add_x_19_3_n136 (.Y(FE_OCPN1908_add_x_19_3_n136), 
	.A(\add_x_19_3/n136 ));
   BUFX4TS FE_OCPC1907_add_x_19_5_n187 (.Y(FE_OCPN1907_add_x_19_5_n187), 
	.A(\add_x_19_5/n187 ));
   CLKBUFX2TS FE_OCPC1906_add_x_19_3_n139 (.Y(FE_OCPN1906_add_x_19_3_n139), 
	.A(\add_x_19_3/n139 ));
   BUFX20TS FE_OCP_DRV_C1894_filesize_29_ (.Y(FE_OCP_DRV_N1894_filesize_29_), 
	.A(filesize[29]));
   CLKBUFX3TS FE_OCPUNCOC1888_n2813 (.Y(FE_OCPUNCON1888_n2813), 
	.A(FE_OCPUNCON1887_n2813));
   BUFX3TS FE_OCPUNCOC1887_n2813 (.Y(FE_OCPUNCON1887_n2813), 
	.A(FE_OCPUNCON1886_n2813));
   BUFX3TS FE_OCPUNCOC1886_n2813 (.Y(FE_OCPUNCON1886_n2813), 
	.A(FE_OCPUNCON1885_n2813));
   BUFX3TS FE_OCPUNCOC1885_n2813 (.Y(FE_OCPUNCON1885_n2813), 
	.A(FE_OCPUNCON1884_n2813));
   BUFX8TS FE_OCPUNCOC1884_n2813 (.Y(FE_OCPUNCON1884_n2813), 
	.A(FE_OCPUNCON1883_n2813));
   BUFX8TS FE_OCPUNCOC1883_n2813 (.Y(FE_OCPUNCON1883_n2813), 
	.A(FE_OCPUNCON1882_n2813));
   BUFX3TS FE_OCPUNCOC1882_n2813 (.Y(FE_OCPUNCON1882_n2813), 
	.A(FE_OCPUNCON1881_n2813));
   BUFX6TS FE_OCPUNCOC1881_n2813 (.Y(FE_OCPUNCON1881_n2813), 
	.A(FE_OCPUNCON1879_n2813));
   BUFX3TS FE_OCPUNCOC1880_n2787 (.Y(FE_OCPUNCON1880_n2787), 
	.A(FE_OCPUNCON1878_n2787));
   BUFX3TS FE_OCPUNCOC1879_n2813 (.Y(FE_OCPUNCON1879_n2813), 
	.A(n2813));
   BUFX3TS FE_OCPUNCOC1878_n2787 (.Y(FE_OCPUNCON1878_n2787), 
	.A(n2787));
   BUFX12TS FE_OCPUNCOC1877_FE_OFN374_offset_22_ (.Y(FE_OCPUNCON1877_FE_OFN374_offset_22_), 
	.A(FE_OFN374_offset_22_));
   BUFX20TS FE_OCPUNCOC1876_offset_22_ (.Y(FE_OCPUNCON1876_offset_22_), 
	.A(offset[22]));
   BUFX20TS FE_OCPUNCOC1875_offset_4_ (.Y(FE_OCPUNCON1875_offset_4_), 
	.A(offset[4]));
   BUFX20TS FE_OCPUNCOC1874_offset_1_ (.Y(FE_OCPUNCON1874_offset_1_), 
	.A(offset[1]));
   BUFX20TS FE_RC_878_0 (.Y(FE_OFN568_offset_28_), 
	.A(offset[28]));
   BUFX20TS FE_RC_877_0 (.Y(FE_OFN410_offset_12_), 
	.A(offset[12]));
   BUFX20TS FE_RC_876_0 (.Y(FE_OFN369_offset_23_), 
	.A(offset[23]));
   BUFX20TS FE_RC_875_0 (.Y(FE_OFN357_offset_26_), 
	.A(offset[26]));
   INVX2TS FE_RC_874_0 (.Y(FE_RN_368_0), 
	.A(\add_x_19_4/n11 ));
   NAND2BX2TS FE_RC_873_0 (.Y(FE_RN_367_0), 
	.B(FE_RN_368_0), 
	.AN(\add_x_19_4/n88 ));
   OAI2BB1X4TS FE_RC_872_0 (.Y(\addr_calc/iir_read_addr[21] ), 
	.B0(FE_RN_367_0), 
	.A1N(\add_x_19_4/n88 ), 
	.A0N(\add_x_19_4/n11 ));
   BUFX20TS FE_OCP_DRV_C1872_filesize_18_ (.Y(FE_OCP_DRV_N1872_filesize_18_), 
	.A(filesize[18]));
   AOI21X2TS FE_RC_853_0 (.Y(\add_x_19_4/n75 ), 
	.B0(\add_x_19_4/n77 ), 
	.A1(\add_x_19_4/n76 ), 
	.A0(\add_x_19_4/n85 ));
   AOI21X4TS FE_RC_851_0 (.Y(\add_x_19_1/n178 ), 
	.B0(\add_x_19_1/n180 ), 
	.A1(\add_x_19_1/n179 ), 
	.A0(\add_x_19_1/n187 ));
   OAI22X4TS FE_RC_845_0 (.Y(\add_x_19_0/n38 ), 
	.B1(n2628), 
	.B0(n1541), 
	.A1(n1541), 
	.A0(\add_x_19_0/n43 ));
   INVX2TS FE_RC_844_0 (.Y(FE_RN_349_0), 
	.A(\add_x_19_0/n36 ));
   NAND2X2TS FE_RC_843_0 (.Y(FE_RN_348_0), 
	.B(FE_RN_349_0), 
	.A(n1541));
   NAND2X2TS FE_RC_842_0 (.Y(FE_RN_347_0), 
	.B(\add_x_19_0/n37 ), 
	.A(FE_RN_348_0));
   NAND2X2TS FE_RC_841_0 (.Y(FE_RN_346_0), 
	.B(\add_x_19_0/n1 ), 
	.A(FE_RN_347_0));
   INVX2TS FE_RC_840_0 (.Y(FE_RN_345_0), 
	.A(\add_x_19_0/n1 ));
   INVX2TS FE_RC_839_0 (.Y(FE_RN_344_0), 
	.A(\add_x_19_0/n36 ));
   OAI21X4TS FE_RC_838_0 (.Y(FE_RN_343_0), 
	.B0(FE_RN_344_0), 
	.A1(n1541), 
	.A0(n2628));
   NAND3X2TS FE_RC_837_0 (.Y(FE_RN_342_0), 
	.C(FE_RN_345_0), 
	.B(\add_x_19_0/n37 ), 
	.A(FE_RN_343_0));
   INVX2TS FE_RC_836_0 (.Y(FE_RN_341_0), 
	.A(\add_x_19_0/n36 ));
   NAND4X4TS FE_RC_835_0 (.Y(FE_RN_340_0), 
	.D(\add_x_19_0/n1 ), 
	.C(FE_RN_341_0), 
	.B(n2628), 
	.A(\add_x_19_0/n43 ));
   INVX2TS FE_RC_834_0 (.Y(FE_RN_339_0), 
	.A(n1541));
   NAND4BBX4TS FE_RC_833_0 (.Y(FE_RN_338_0), 
	.D(FE_RN_339_0), 
	.C(\add_x_19_0/n37 ), 
	.BN(\add_x_19_0/n1 ), 
	.AN(\add_x_19_0/n43 ));
   NAND4X4TS FE_RC_832_0 (.Y(\addr_calc/fft_read_addr[31] ), 
	.D(FE_RN_346_0), 
	.C(FE_RN_342_0), 
	.B(FE_RN_340_0), 
	.A(FE_RN_338_0));
   BUFX20TS FE_RC_791_0 (.Y(FE_OFN422_offset_9_), 
	.A(offset[9]));
   BUFX20TS FE_RC_790_0 (.Y(FE_OFN424_offset_9_), 
	.A(offset[9]));
   NOR2X8TS FE_RC_789_0 (.Y(\add_x_19_5/n151 ), 
	.B(\addr_calc/iir_write_calc/count[9] ), 
	.A(offset[9]));
   BUFX20TS FE_RC_786_0 (.Y(FE_OCP_RBN1842_offset_7_), 
	.A(offset[7]));
   BUFX20TS FE_OCP_RBC1841_offset_7_ (.Y(FE_OCP_RBN1841_offset_7_), 
	.A(FE_OCP_RBN1842_offset_7_));
   BUFX20TS FE_OCP_RBC1840_offset_7_ (.Y(FE_OCP_RBN1840_offset_7_), 
	.A(FE_OCP_RBN1842_offset_7_));
   CLKBUFX2TS FE_OCPC1825_add_x_19_3_n68 (.Y(FE_OCPN1825_add_x_19_3_n68), 
	.A(\add_x_19_3/n68 ));
   BUFX20TS FE_OCP_DRV_C1824_filesize_19_ (.Y(FE_OCP_DRV_N1824_filesize_19_), 
	.A(filesize[19]));
   BUFX20TS FE_OCP_DRV_C1818_filesize_20_ (.Y(FE_OCP_DRV_N1818_filesize_20_), 
	.A(filesize[20]));
   NAND2X2TS FE_RC_780_0 (.Y(FE_RN_310_0), 
	.B(n1229), 
	.A(\add_x_19_2/n60 ));
   NAND2X2TS FE_RC_779_0 (.Y(n1228), 
	.B(n1230), 
	.A(FE_RN_310_0));
   OAI21X4TS FE_RC_776_0 (.Y(\add_x_19_5/n157 ), 
	.B0(FE_RN_104_0), 
	.A1(FE_RN_107_0), 
	.A0(FE_RN_106_0));
   OAI21X2TS FE_RC_771_0 (.Y(n1548), 
	.B0(\add_x_19_2/n182 ), 
	.A1(\add_x_19_2/n181 ), 
	.A0(\add_x_19_2/n185 ));
   CLKINVX4TS FE_OCP_RBC1788_add_x_19_3_n163 (.Y(FE_OCP_RBN1788_add_x_19_3_n163), 
	.A(FE_OCP_RBN1787_add_x_19_3_n163));
   CLKBUFX2TS FE_OCP_RBC1787_add_x_19_3_n163 (.Y(FE_OCP_RBN1787_add_x_19_3_n163), 
	.A(\add_x_19_3/n163 ));
   CLKBUFX3TS FE_OCPUNCOC1750_offset_1_ (.Y(FE_OCPUNCON1750_offset_1_), 
	.A(offset[1]));
   BUFX20TS FE_RC_765_0 (.Y(FE_OFN353_offset_27_), 
	.A(offset[27]));
   BUFX8TS FE_OCPC1732_n1718 (.Y(FE_OCPN1732_n1718), 
	.A(n1718));
   BUFX16TS FE_OCPC1731_FE_OCPUNCON1650_add_x_19_4_n43 (.Y(FE_OCPN1731_FE_OCPUNCON1650_add_x_19_4_n43), 
	.A(FE_OCPUNCON1650_add_x_19_4_n43));
   BUFX3TS FE_OCPC1730_add_x_19_0_n43 (.Y(FE_OCPN1730_add_x_19_0_n43), 
	.A(\add_x_19_0/n43 ));
   BUFX3TS FE_OCPC1729_FE_OFN528_add_x_19_0_n113 (.Y(FE_OCPN1729_FE_OFN528_add_x_19_0_n113), 
	.A(FE_OCPN1728_FE_OFN528_add_x_19_0_n113));
   BUFX12TS FE_OCPC1728_FE_OFN528_add_x_19_0_n113 (.Y(FE_OCPN1728_FE_OFN528_add_x_19_0_n113), 
	.A(FE_OFN528_add_x_19_0_n113));
   BUFX20TS FE_OCPUNCOC1686_offset_20_ (.Y(FE_OCPUNCON1686_offset_20_), 
	.A(offset[20]));
   NAND2X6TS FE_RC_764_0 (.Y(FE_OFN541_addr_calc_iir_read_addr_9_), 
	.B(FE_RN_188_0), 
	.A(FE_RN_269_0));
   XNOR2X4TS FE_RC_763_0 (.Y(FE_OFN118_addr_calc_iir_read_addr_15_), 
	.B(\add_x_19_4/n17 ), 
	.A(\add_x_19_4/n122 ));
   BUFX20TS FE_RC_758_0 (.Y(FE_OFN614_filesize_1_), 
	.A(filesize[1]));
   BUFX20TS FE_RC_757_0 (.Y(FE_OFN613_filesize_2_), 
	.A(filesize[2]));
   BUFX20TS FE_RC_756_0 (.Y(FE_OFN580_offset_16_), 
	.A(offset[16]));
   BUFX20TS FE_RC_751_0 (.Y(FE_OFN386_offset_18_), 
	.A(offset[18]));
   BUFX20TS FE_RC_749_0 (.Y(FE_OFN365_offset_24_), 
	.A(offset[24]));
   BUFX20TS FE_RC_748_0 (.Y(FE_OFN361_offset_25_), 
	.A(offset[25]));
   NOR2X2TS FE_RC_744_0 (.Y(FE_RN_304_0), 
	.B(n1567), 
	.A(\add_x_19_4/n135 ));
   OAI21X2TS FE_RC_743_0 (.Y(FE_RN_303_0), 
	.B0(\add_x_19_4/n121 ), 
	.A1(\add_x_19_4/n120 ), 
	.A0(\add_x_19_4/n124 ));
   AOI21X1TS FE_RC_742_0 (.Y(FE_RN_302_0), 
	.B0(FE_RN_303_0), 
	.A1(\add_x_19_4/n127 ), 
	.A0(n1549));
   OAI21X2TS FE_RC_741_0 (.Y(FE_RN_301_0), 
	.B0(FE_RN_302_0), 
	.A1(n1567), 
	.A0(\add_x_19_4/n136 ));
   AOI21X4TS FE_RC_740_0 (.Y(\add_x_19_4/n113 ), 
	.B0(FE_RN_301_0), 
	.A1(FE_RN_304_0), 
	.A0(FE_OCP_RBN1981_add_x_19_4_n157));
   OAI21X4TS FE_RC_727_0 (.Y(\add_x_19_5/n104 ), 
	.B0(\add_x_19_5/n106 ), 
	.A1(\add_x_19_5/n105 ), 
	.A0(\add_x_19_5/n111 ));
   NOR3BX1TS FE_RC_725_0 (.Y(FE_RN_294_0), 
	.C(\add_x_19_4/n40 ), 
	.B(n2634), 
	.AN(n1640));
   AOI2BB1X1TS FE_RC_724_0 (.Y(FE_RN_293_0), 
	.B0(FE_RN_294_0), 
	.A1N(n1583), 
	.A0N(n1640));
   NOR2BX1TS FE_RC_723_0 (.Y(FE_RN_292_0), 
	.B(n1640), 
	.AN(n2634));
   NAND2X4TS FE_RC_722_0 (.Y(FE_RN_291_0), 
	.B(FE_RN_292_0), 
	.A(FE_OCPN1731_FE_OCPUNCON1650_add_x_19_4_n43));
   AND2X2TS FE_RC_721_0 (.Y(FE_RN_290_0), 
	.B(n1583), 
	.A(n1640));
   NAND2BX4TS FE_RC_720_0 (.Y(FE_RN_289_0), 
	.B(FE_RN_290_0), 
	.AN(FE_OCPN1731_FE_OCPUNCON1650_add_x_19_4_n43));
   NAND3X6TS FE_RC_719_0 (.Y(\addr_calc/iir_read_addr[30] ), 
	.C(FE_RN_293_0), 
	.B(FE_RN_291_0), 
	.A(FE_RN_289_0));
   INVX2TS FE_RC_714_0 (.Y(FE_RN_285_0), 
	.A(\add_x_19_3/n72 ));
   NOR2X4TS FE_RC_713_0 (.Y(FE_RN_284_0), 
	.B(FE_RN_285_0), 
	.A(\add_x_19_3/n113 ));
   OR2X8TS FE_RC_712_0 (.Y(\add_x_19_3/n69 ), 
	.B(\add_x_19_3/n73 ), 
	.A(FE_RN_284_0));
   NAND2X2TS FE_RC_692_0 (.Y(FE_RN_269_0), 
	.B(FE_RN_208_0), 
	.A(FE_RN_207_0));
   OAI21X4TS FE_RC_689_0 (.Y(\add_x_19_4/n43 ), 
	.B0(\add_x_19_4/n45 ), 
	.A1(\add_x_19_4/n44 ), 
	.A0(FE_OFN527_add_x_19_4_n113));
   OAI21X4TS FE_RC_688_0 (.Y(\add_x_19_4/n157 ), 
	.B0(\add_x_19_4/n159 ), 
	.A1(\add_x_19_4/n158 ), 
	.A0(\add_x_19_4/n178 ));
   NAND2X6TS FE_RC_646_0 (.Y(n2589), 
	.B(\DP_OP_158_296_6262/n1986 ), 
	.A(\DP_OP_158_296_6262/n1931 ));
   NAND2X8TS FE_RC_645_0 (.Y(FE_OCPUNCON1081_n2589), 
	.B(\DP_OP_158_296_6262/n1931 ), 
	.A(\DP_OP_158_296_6262/n1986 ));
   INVX2TS FE_RC_638_0 (.Y(FE_RN_241_0), 
	.A(\add_x_19_4/n219 ));
   OAI21X4TS FE_RC_637_0 (.Y(n1397), 
	.B0(\add_x_19_4/n176 ), 
	.A1(FE_RN_241_0), 
	.A0(FE_OCP_RBN1979_add_x_19_4_n178));
   INVX2TS FE_RC_636_0 (.Y(FE_RN_240_0), 
	.A(\add_x_19_4/n170 ));
   NAND2BX2TS FE_RC_635_0 (.Y(FE_RN_239_0), 
	.B(FE_RN_240_0), 
	.AN(n1398));
   INVX2TS FE_RC_634_0 (.Y(FE_RN_238_0), 
	.A(\add_x_19_4/n219 ));
   AOI22X2TS FE_RC_633_0 (.Y(FE_RN_237_0), 
	.B1(FE_RN_238_0), 
	.B0(\add_x_19_4/n176 ), 
	.A1(\add_x_19_4/n176 ), 
	.A0(FE_OCP_RBN1979_add_x_19_4_n178));
   NAND2X2TS FE_RC_632_0 (.Y(n1399), 
	.B(FE_RN_239_0), 
	.A(FE_RN_237_0));
   CLKINVX4TS FE_RC_601_0 (.Y(\add_x_19_0/n66 ), 
	.A(FE_RN_217_0));
   INVX2TS FE_RC_600_0 (.Y(FE_RN_219_0), 
	.A(\add_x_19_0/n63 ));
   INVX2TS FE_RC_599_0 (.Y(FE_RN_218_0), 
	.A(n2038));
   NAND2BX4TS FE_RC_598_0 (.Y(FE_RN_217_0), 
	.B(FE_RN_218_0), 
	.AN(FE_OFN368_offset_24_));
   AND2X6TS FE_RC_597_0 (.Y(\add_x_19_0/n61 ), 
	.B(FE_RN_219_0), 
	.A(FE_RN_217_0));
   NAND2X8TS FE_RC_590_0 (.Y(\add_x_19_1/n176 ), 
	.B(\addr_calc/fft_write_calc/count[4] ), 
	.A(offset[4]));
   INVX2TS FE_RC_589_0 (.Y(FE_RN_214_0), 
	.A(offset[4]));
   INVX2TS FE_RC_588_0 (.Y(FE_RN_213_0), 
	.A(\addr_calc/fft_write_calc/count[4] ));
   OAI31X2TS FE_RC_587_0 (.Y(\add_x_19_1/n169 ), 
	.B0(\add_x_19_1/n171 ), 
	.A2(FE_RN_213_0), 
	.A1(FE_RN_214_0), 
	.A0(\add_x_19_1/n170 ));
   BUFX20TS FE_RC_586_0 (.Y(FE_OCPUNCON1564_offset_5_), 
	.A(offset[5]));
   NOR2X8TS FE_RC_585_0 (.Y(\add_x_19_2/n170 ), 
	.B(offset[5]), 
	.A(\addr_calc/fir_read_calc/count[5] ));
   BUFX16TS FE_OCPUNCOC1650_add_x_19_4_n43 (.Y(FE_OCPUNCON1650_add_x_19_4_n43), 
	.A(\add_x_19_4/n43 ));
   INVX8TS FE_RC_583_0 (.Y(n2602), 
	.A(FE_RN_212_0));
   XNOR2X4TS FE_RC_582_0 (.Y(FE_RN_212_0), 
	.B(n1678), 
	.A(n1736));
   CLKINVX2TS FE_RC_575_0 (.Y(FE_RN_208_0), 
	.A(FE_RN_86_0));
   INVX2TS FE_RC_574_0 (.Y(FE_RN_207_0), 
	.A(n1409));
   OAI21X2TS FE_RC_572_0 (.Y(\add_x_19_2/n99 ), 
	.B0(\add_x_19_2/n101 ), 
	.A1(\add_x_19_2/n100 ), 
	.A0(\add_x_19_2/n102 ));
   XOR2X4TS FE_RC_571_0 (.Y(\addr_calc/fir_read_addr[17] ), 
	.B(\add_x_19_2/n15 ), 
	.A(\add_x_19_2/n107 ));
   XOR2X4TS FE_RC_569_0 (.Y(\addr_calc/fft_write_addr[20] ), 
	.B(n1441), 
	.A(\add_x_19_1/n91 ));
   XOR2X4TS FE_RC_567_0 (.Y(\addr_calc/fft_write_addr[17] ), 
	.B(n1385), 
	.A(n1384));
   OAI21X4TS FE_RC_566_0 (.Y(n1568), 
	.B0(\add_x_19_2/n90 ), 
	.A1(\add_x_19_2/n89 ), 
	.A0(\add_x_19_2/n91 ));
   AOI21X4TS FE_RC_564_0 (.Y(\add_x_19_4/n107 ), 
	.B0(\add_x_19_4/n109 ), 
	.A1(\add_x_19_4/n207 ), 
	.A0(\add_x_19_4/n112 ));
   OAI21X4TS FE_RC_562_0 (.Y(\add_x_19_0/n130 ), 
	.B0(\add_x_19_0/n132 ), 
	.A1(\add_x_19_0/n131 ), 
	.A0(\add_x_19_0/n133 ));
   NAND3X8TS FE_RC_551_0 (.Y(FE_OFN525_add_x_19_3_n157), 
	.C(FE_RN_108_0), 
	.B(FE_RN_109_0), 
	.A(FE_RN_111_0));
   NAND3X4TS FE_RC_550_0 (.Y(FE_RN_100_0), 
	.C(n1558), 
	.B(\add_x_19_0/n168 ), 
	.A(FE_RN_101_0));
   NAND3X6TS FE_RC_549_0 (.Y(FE_RN_109_0), 
	.C(\add_x_19_3/n160 ), 
	.B(\add_x_19_3/n168 ), 
	.A(FE_RN_110_0));
   OAI21X4TS FE_RC_546_0 (.Y(\add_x_19_1/n157 ), 
	.B0(\add_x_19_1/n159 ), 
	.A1(\add_x_19_1/n158 ), 
	.A0(\add_x_19_1/n178 ));
   AOI21X4TS FE_RC_545_0 (.Y(FE_RN_106_0), 
	.B0(\add_x_19_5/n180 ), 
	.A1(\add_x_19_5/n187 ), 
	.A0(\add_x_19_5/n179 ));
   CLKBUFX3TS FE_OCPUNCOC1576_n2812 (.Y(FE_OCPUNCON1576_n2812), 
	.A(FE_OCPUNCON1575_n2812));
   BUFX4TS FE_OCPUNCOC1575_n2812 (.Y(FE_OCPUNCON1575_n2812), 
	.A(FE_OCPUNCON1574_n2812));
   BUFX2TS FE_OCPUNCOC1574_n2812 (.Y(FE_OCPUNCON1574_n2812), 
	.A(FE_OCPUNCON1573_n2812));
   BUFX4TS FE_OCPUNCOC1573_n2812 (.Y(FE_OCPUNCON1573_n2812), 
	.A(FE_OCPUNCON1572_n2812));
   BUFX3TS FE_OCPUNCOC1572_n2812 (.Y(FE_OCPUNCON1572_n2812), 
	.A(FE_OCPUNCON1571_n2812));
   BUFX3TS FE_OCPUNCOC1571_n2812 (.Y(FE_OCPUNCON1571_n2812), 
	.A(FE_OCPUNCON1570_n2812));
   BUFX4TS FE_OCPUNCOC1570_n2812 (.Y(FE_OCPUNCON1570_n2812), 
	.A(FE_OCPUNCON1569_n2812));
   BUFX6TS FE_OCPUNCOC1569_n2812 (.Y(FE_OCPUNCON1569_n2812), 
	.A(FE_OCPUNCON1568_n2812));
   BUFX3TS FE_OCPUNCOC1568_n2812 (.Y(FE_OCPUNCON1568_n2812), 
	.A(n2812));
   BUFX8TS FE_OCPUNCOC1567_n1717 (.Y(FE_OCPUNCON1567_n1717), 
	.A(n1717));
   CLKBUFX2TS FE_OCPUNCOC1562_filesize_10_ (.Y(FE_OCPUNCON1562_filesize_10_), 
	.A(filesize[10]));
   AND2X8TS FE_RC_541_0 (.Y(n787), 
	.B(n1780), 
	.A(n1779));
   XNOR2X4TS FE_RC_540_0 (.Y(FE_OFN126_addr_calc_iir_write_addr_25_), 
	.B(\add_x_19_5/n7 ), 
	.A(\add_x_19_5/n65 ));
   XNOR2X4TS FE_RC_538_0 (.Y(FE_OFN116_addr_calc_iir_read_addr_24_), 
	.B(n1467), 
	.A(n1611));
   OA21X4TS FE_RC_537_0 (.Y(\add_x_19_0/n133 ), 
	.B0(\add_x_19_0/n136 ), 
	.A1(\add_x_19_0/n135 ), 
	.A0(\add_x_19_0/n156 ));
   BUFX20TS FE_RC_535_0 (.Y(FE_OFN481_filesize_16_), 
	.A(FE_OCP_DRV_N1389_filesize_16_));
   BUFX20TS FE_RC_531_0 (.Y(FE_OCPUNCON1062_offset_19_), 
	.A(offset[19]));
   NAND2X2TS FE_RC_526_0 (.Y(FE_RN_205_0), 
	.B(\add_x_19_5/n9 ), 
	.A(\add_x_19_5/n80 ));
   NAND2X6TS FE_RC_525_0 (.Y(\addr_calc/iir_write_addr[23] ), 
	.B(FE_RN_205_0), 
	.A(FE_RN_161_0));
   CLKINVX12TS FE_RC_522_0 (.Y(n1778), 
	.A(FE_RN_203_0));
   XOR2X4TS FE_RC_521_0 (.Y(FE_RN_203_0), 
	.B(n2325), 
	.A(\DP_OP_158_296_6262/n1826 ));
   OAI21X4TS FE_RC_520_0 (.Y(\add_x_19_0/n65 ), 
	.B0(\add_x_19_0/n67 ), 
	.A1(\add_x_19_0/n66 ), 
	.A0(\add_x_19_0/n68 ));
   XOR2X4TS FE_RC_519_0 (.Y(n1564), 
	.B(\addr_calc/iir_write_calc/count[30] ), 
	.A(n2625));
   INVX2TS FE_RC_518_0 (.Y(FE_RN_202_0), 
	.A(\add_x_19_3/n128 ));
   CLKINVX1TS FE_RC_517_0 (.Y(FE_RN_201_0), 
	.A(n1301));
   OAI2BB1X1TS FE_RC_516_0 (.Y(n1302), 
	.B0(n1300), 
	.A1N(FE_RN_201_0), 
	.A0N(FE_RN_202_0));
   XOR2X4TS FE_RC_515_0 (.Y(\addr_calc/iir_write_addr[30] ), 
	.B(n1359), 
	.A(n1358));
   INVX2TS FE_RC_514_0 (.Y(FE_RN_200_0), 
	.A(\add_x_19_1/n7 ));
   NAND2BX2TS FE_RC_513_0 (.Y(FE_RN_199_0), 
	.B(FE_RN_200_0), 
	.AN(\add_x_19_1/n65 ));
   OAI2BB1X4TS FE_RC_512_0 (.Y(\addr_calc/fft_write_addr[25] ), 
	.B0(FE_RN_199_0), 
	.A1N(\add_x_19_1/n65 ), 
	.A0N(\add_x_19_1/n7 ));
   INVX2TS FE_RC_511_0 (.Y(FE_RN_198_0), 
	.A(\add_x_19_1/n4 ));
   NAND2BX2TS FE_RC_510_0 (.Y(FE_RN_197_0), 
	.B(FE_RN_198_0), 
	.AN(\add_x_19_1/n50 ));
   OAI2BB1X4TS FE_RC_509_0 (.Y(\addr_calc/fft_write_addr[28] ), 
	.B0(FE_RN_197_0), 
	.A1N(\add_x_19_1/n50 ), 
	.A0N(\add_x_19_1/n4 ));
   OAI21X2TS FE_RC_504_0 (.Y(\add_x_19_3/n35 ), 
	.B0(\add_x_19_3/n37 ), 
	.A1(\add_x_19_3/n36 ), 
	.A0(\add_x_19_3/n38 ));
   NAND2X2TS FE_RC_497_0 (.Y(FE_RN_192_0), 
	.B(n1552), 
	.A(\add_x_19_1/n38 ));
   NAND2X2TS FE_RC_496_0 (.Y(n1551), 
	.B(n1553), 
	.A(FE_RN_192_0));
   XOR2X4TS FE_RC_495_0 (.Y(\addr_calc/fir_read_addr[20] ), 
	.B(n1404), 
	.A(\add_x_19_2/n91 ));
   OR2X2TS FE_RC_494_0 (.Y(FE_RN_191_0), 
	.B(\add_x_19_0/n151 ), 
	.A(n1418));
   NOR2X2TS FE_RC_493_0 (.Y(FE_RN_190_0), 
	.B(FE_RN_191_0), 
	.A(n1417));
   NAND2BX4TS FE_RC_492_0 (.Y(\addr_calc/fft_read_addr[9] ), 
	.B(n1419), 
	.AN(FE_RN_190_0));
   XOR2X4TS FE_RC_491_0 (.Y(\addr_calc/fir_write_addr[20] ), 
	.B(n1438), 
	.A(FE_OCP_RBN1381_add_x_19_3_n92));
   NAND2X2TS FE_RC_488_0 (.Y(FE_RN_188_0), 
	.B(FE_RN_87_0), 
	.A(n1409));
   OAI21X2TS FE_RC_486_0 (.Y(\add_x_19_2/n130 ), 
	.B0(\add_x_19_2/n132 ), 
	.A1(\add_x_19_2/n131 ), 
	.A0(\add_x_19_2/n133 ));
   AOI21X4TS FE_RC_485_0 (.Y(\add_x_19_1/n102 ), 
	.B0(\add_x_19_1/n104 ), 
	.A1(\add_x_19_1/n103 ), 
	.A0(\add_x_19_1/n112 ));
   XOR2X4TS FE_RC_484_0 (.Y(\addr_calc/fir_read_addr[12] ), 
	.B(n1363), 
	.A(\add_x_19_2/n133 ));
   OAI21X4TS FE_RC_472_0 (.Y(\add_x_19_4/n134 ), 
	.B0(\add_x_19_4/n136 ), 
	.A1(\add_x_19_4/n135 ), 
	.A0(FE_OCP_RBN1925_add_x_19_4_n157));
   AOI21X2TS FE_RC_470_0 (.Y(\add_x_19_4/n45 ), 
	.B0(\add_x_19_4/n47 ), 
	.A1(\add_x_19_4/n46 ), 
	.A0(\add_x_19_4/n73 ));
   OAI21X2TS FE_RC_468_0 (.Y(\add_x_19_1/n73 ), 
	.B0(FE_RN_152_0), 
	.A1(\add_x_19_1/n74 ), 
	.A0(\add_x_19_1/n94 ));
   AOI21X4TS FE_RC_466_0 (.Y(\add_x_19_0/n94 ), 
	.B0(FE_RN_64_0), 
	.A1(\add_x_19_0/n104 ), 
	.A0(\add_x_19_0/n95 ));
   OAI21X4TS FE_RC_463_0 (.Y(\add_x_19_4/n104 ), 
	.B0(\add_x_19_4/n106 ), 
	.A1(\add_x_19_4/n105 ), 
	.A0(\add_x_19_4/n111 ));
   AOI21X4TS FE_RC_460_0 (.Y(\add_x_19_2/n52 ), 
	.B0(\add_x_19_2/n54 ), 
	.A1(\add_x_19_2/n53 ), 
	.A0(\add_x_19_2/n62 ));
   AOI21X4TS FE_RC_459_0 (.Y(n1594), 
	.B0(n1595), 
	.A1(\add_x_19_3/n118 ), 
	.A0(\add_x_19_3/n127 ));
   CLKINVX6TS FE_RC_458_0 (.Y(FE_RN_111_0), 
	.A(FE_RN_187_0));
   OAI21X2TS FE_RC_457_0 (.Y(FE_RN_187_0), 
	.B0(\add_x_19_3/n163 ), 
	.A1(\add_x_19_3/n166 ), 
	.A0(\add_x_19_3/n162 ));
   AOI21X4TS FE_RC_456_0 (.Y(FE_RN_104_0), 
	.B0(FE_RN_105_0), 
	.A1(\add_x_19_5/n169 ), 
	.A0(\add_x_19_5/n160 ));
   OAI21X2TS FE_RC_454_0 (.Y(\add_x_19_2/n104 ), 
	.B0(\add_x_19_2/n106 ), 
	.A1(\add_x_19_2/n105 ), 
	.A0(\add_x_19_2/n111 ));
   OAI21X2TS FE_RC_453_0 (.Y(\add_x_19_5/n180 ), 
	.B0(\add_x_19_5/n182 ), 
	.A1(\add_x_19_5/n185 ), 
	.A0(\add_x_19_5/n181 ));
   BUFX6TS FE_OCP_RBC1495_offset_5_ (.Y(FE_OCP_RBN1495_offset_5_), 
	.A(FE_OCPUNCON1564_offset_5_));
   BUFX8TS FE_OCP_RBC1494_offset_5_ (.Y(FE_OCP_RBN1494_offset_5_), 
	.A(FE_OCPUNCON1564_offset_5_));
   BUFX16TS FE_OCP_RBC1493_offset_5_ (.Y(FE_OCP_RBN1493_offset_5_), 
	.A(FE_OCP_RBN1494_offset_5_));
   BUFX20TS FE_OCP_RBC1492_offset_5_ (.Y(FE_OCP_RBN1492_offset_5_), 
	.A(FE_OCP_RBN1494_offset_5_));
   BUFX16TS FE_OCPUNCOC1425_FE_OFN443_offset_4_ (.Y(FE_OCPUNCON1425_FE_OFN443_offset_4_), 
	.A(FE_OFN443_offset_4_));
   BUFX20TS FE_OCP_DRV_C1389_filesize_16_ (.Y(FE_OCP_DRV_N1389_filesize_16_), 
	.A(filesize[16]));
   AOI21X4TS FE_RC_440_0 (.Y(n1384), 
	.B0(\add_x_19_1/n109 ), 
	.A1(\add_x_19_1/n207 ), 
	.A0(\add_x_19_1/n112 ));
   OAI21X4TS FE_RC_439_0 (.Y(\add_x_19_4/n146 ), 
	.B0(\add_x_19_4/n148 ), 
	.A1(\add_x_19_4/n147 ), 
	.A0(FE_OCP_RBN1925_add_x_19_4_n157));
   AOI21X4TS FE_RC_436_0 (.Y(n1299), 
	.B0(\add_x_19_3/n47 ), 
	.A1(\add_x_19_3/n46 ), 
	.A0(\add_x_19_3/n73 ));
   OAI21X2TS FE_RC_425_0 (.Y(\add_x_19_2/n54 ), 
	.B0(\add_x_19_2/n56 ), 
	.A1(FE_OFN142_add_x_19_2_n59), 
	.A0(\add_x_19_2/n55 ));
   CLKINVX6TS FE_OCP_RBC1383_add_x_19_0_n92 (.Y(FE_OCP_RBN1383_add_x_19_0_n92), 
	.A(\add_x_19_0/n92 ));
   INVX3TS FE_OCP_RBC1381_add_x_19_3_n92 (.Y(FE_OCP_RBN1381_add_x_19_3_n92), 
	.A(\add_x_19_3/n92 ));
   CLKINVX6TS FE_OCP_RBC1379_add_x_19_1_n69 (.Y(FE_OCP_RBN1379_add_x_19_1_n69), 
	.A(\add_x_19_1/n69 ));
   INVX6TS FE_OCP_RBC1378_add_x_19_3_n113 (.Y(FE_OCP_RBN1378_add_x_19_3_n113), 
	.A(\add_x_19_3/n113 ));
   CLKINVX12TS FE_OCP_RBC1366_FE_OCP_DRV_N1167_offset_20_ (.Y(FE_OCP_RBN1366_FE_OCP_DRV_N1167_offset_20_), 
	.A(FE_OCPUNCON1686_offset_20_));
   CLKINVX1TS FE_OCP_RBC1365_FE_OCP_DRV_N1167_offset_20_ (.Y(FE_OCP_RBN1365_FE_OCP_DRV_N1167_offset_20_), 
	.A(FE_OCPUNCON1686_offset_20_));
   CLKINVX12TS FE_OCP_RBC1364_FE_OCP_DRV_N1167_offset_20_ (.Y(FE_OCP_RBN1364_FE_OCP_DRV_N1167_offset_20_), 
	.A(FE_OCPUNCON1686_offset_20_));
   CLKINVX2TS FE_OCP_RBC1363_FE_OCP_DRV_N1167_offset_20_ (.Y(FE_OCP_RBN1363_FE_OCP_DRV_N1167_offset_20_), 
	.A(FE_OCPUNCON1686_offset_20_));
   BUFX3TS FE_OCPC1362_add_x_19_2_n83 (.Y(FE_OCPN1362_add_x_19_2_n83), 
	.A(\add_x_19_2/n83 ));
   BUFX20TS FE_OCP_DRV_C1336_filesize_0_ (.Y(FE_OCP_DRV_N1336_filesize_0_), 
	.A(filesize[0]));
   BUFX3TS FE_OCPUNCOC1318_FE_OFN361_offset_25_ (.Y(FE_OCPUNCON1318_FE_OFN361_offset_25_), 
	.A(FE_OFN361_offset_25_));
   BUFX20TS FE_OCPUNCOC1278_offset_7_ (.Y(FE_OCPUNCON1278_offset_7_), 
	.A(FE_OCP_RBN1841_offset_7_));
   CLKBUFX2TS FE_OCPC1257_add_x_19_0_n162 (.Y(FE_OCPN1257_add_x_19_0_n162), 
	.A(\add_x_19_0/n162 ));
   CLKBUFX2TS FE_OCPC1256_add_x_19_3_n162 (.Y(FE_OCPN1256_add_x_19_3_n162), 
	.A(\add_x_19_3/n162 ));
   CLKBUFX2TS FE_OCPC1255_add_x_19_3_n181 (.Y(FE_OCPN1255_add_x_19_3_n181), 
	.A(\add_x_19_3/n181 ));
   BUFX8TS FE_OCPC1230_n1611 (.Y(FE_OCPN1230_n1611), 
	.A(n1611));
   BUFX8TS FE_OCPC1229_add_x_19_5_n68 (.Y(FE_OCPN1229_add_x_19_5_n68), 
	.A(\add_x_19_5/n68 ));
   BUFX3TS FE_OCPC1226_add_x_19_4_n112 (.Y(FE_OCPN1226_add_x_19_4_n112), 
	.A(\add_x_19_4/n112 ));
   CLKBUFX2TS FE_OCPC1225_add_x_19_5_n170 (.Y(FE_OCPN1225_add_x_19_5_n170), 
	.A(\add_x_19_5/n170 ));
   BUFX4TS FE_OCPC1224_FE_OFN445_offset_4_ (.Y(FE_OCPN1224_FE_OFN445_offset_4_), 
	.A(FE_OCPUNCON1425_FE_OFN443_offset_4_));
   CLKBUFX2TS FE_OCPC1223_add_x_19_1_n181 (.Y(FE_OCPN1223_add_x_19_1_n181), 
	.A(\add_x_19_1/n181 ));
   CLKBUFX2TS FE_OCPC1222_add_x_19_5_n162 (.Y(FE_OCPN1222_add_x_19_5_n162), 
	.A(\add_x_19_5/n162 ));
   CLKBUFX2TS FE_OCPC1221_add_x_19_4_n162 (.Y(FE_OCPN1221_add_x_19_4_n162), 
	.A(\add_x_19_4/n162 ));
   CLKBUFX2TS FE_OCPC1220_add_x_19_2_n181 (.Y(FE_OCPN1220_add_x_19_2_n181), 
	.A(\add_x_19_2/n181 ));
   CLKBUFX2TS FE_OCPC1189_add_x_19_0_n181 (.Y(FE_OCPN1189_add_x_19_0_n181), 
	.A(\add_x_19_0/n181 ));
   BUFX16TS FE_OCPC1188_offset_3_ (.Y(FE_OCPN1188_offset_3_), 
	.A(FE_OCPUNCON1563_offset_3_));
   BUFX20TS FE_OCP_DRV_C1099_filesize_14_ (.Y(FE_OCP_DRV_N1099_filesize_14_), 
	.A(filesize[14]));
   BUFX3TS FE_OCPUNCOC1093_n2805 (.Y(FE_OCPUNCON1093_n2805), 
	.A(FE_OCPUNCON1092_n2805));
   BUFX3TS FE_OCPUNCOC1092_n2805 (.Y(FE_OCPUNCON1092_n2805), 
	.A(FE_OCPUNCON1091_n2805));
   BUFX3TS FE_OCPUNCOC1091_n2805 (.Y(FE_OCPUNCON1091_n2805), 
	.A(FE_OCPUNCON1090_n2805));
   BUFX3TS FE_OCPUNCOC1090_n2805 (.Y(FE_OCPUNCON1090_n2805), 
	.A(FE_OCPUNCON1089_n2805));
   BUFX3TS FE_OCPUNCOC1089_n2805 (.Y(FE_OCPUNCON1089_n2805), 
	.A(FE_OCPUNCON1088_n2805));
   BUFX8TS FE_OCPUNCOC1088_n2805 (.Y(FE_OCPUNCON1088_n2805), 
	.A(FE_OCPUNCON1087_n2805));
   BUFX3TS FE_OCPUNCOC1087_n2805 (.Y(FE_OCPUNCON1087_n2805), 
	.A(FE_OCPUNCON1086_n2805));
   BUFX3TS FE_OCPUNCOC1086_n2805 (.Y(FE_OCPUNCON1086_n2805), 
	.A(FE_OCPUNCON1085_n2805));
   BUFX3TS FE_OCPUNCOC1085_n2805 (.Y(FE_OCPUNCON1085_n2805), 
	.A(FE_OCPUNCON1084_n2805));
   BUFX3TS FE_OCPUNCOC1084_n2805 (.Y(FE_OCPUNCON1084_n2805), 
	.A(FE_OCPUNCON1083_n2805));
   BUFX3TS FE_OCPUNCOC1083_n2805 (.Y(FE_OCPUNCON1083_n2805), 
	.A(n2805));
   BUFX16TS FE_OCPUNCOC1082_n2589 (.Y(FE_OCPUNCON1082_n2589), 
	.A(FE_OCPUNCON1081_n2589));
   BUFX12TS FE_OCPUNCOC1080_FE_OFN386_offset_18_ (.Y(FE_OCPUNCON1080_FE_OFN386_offset_18_), 
	.A(FE_OCPUNCON1072_FE_OFN386_offset_18_));
   BUFX8TS FE_OCPUNCOC1079_FE_OFN382_offset_19_ (.Y(FE_OCPUNCON1079_FE_OFN382_offset_19_), 
	.A(FE_OCPUNCON1071_FE_OFN382_offset_19_));
   BUFX8TS FE_OCPUNCOC1078_FE_OFN377_offset_21_ (.Y(FE_OCPUNCON1078_FE_OFN377_offset_21_), 
	.A(FE_OCPUNCON1070_FE_OFN377_offset_21_));
   BUFX16TS FE_OCPUNCOC1077_FE_OFN459_offset_0_ (.Y(FE_OCPUNCON1077_FE_OFN459_offset_0_), 
	.A(FE_OFN459_offset_0_));
   BUFX16TS FE_OCPUNCOC1076_FE_OFN451_offset_2_ (.Y(FE_OCPUNCON1076_FE_OFN451_offset_2_), 
	.A(FE_OFN451_offset_2_));
   BUFX20TS FE_OCPUNCOC1075_FE_OFN447_offset_3_ (.Y(FE_OCPUNCON1075_FE_OFN447_offset_3_), 
	.A(FE_OFN447_offset_3_));
   BUFX16TS FE_OCPUNCOC1073_FE_OFN410_offset_12_ (.Y(FE_OCPUNCON1073_FE_OFN410_offset_12_), 
	.A(FE_OFN410_offset_12_));
   BUFX4TS FE_OCPUNCOC1072_FE_OFN386_offset_18_ (.Y(FE_OCPUNCON1072_FE_OFN386_offset_18_), 
	.A(FE_OFN386_offset_18_));
   BUFX3TS FE_OCPUNCOC1071_FE_OFN382_offset_19_ (.Y(FE_OCPUNCON1071_FE_OFN382_offset_19_), 
	.A(FE_OFN382_offset_19_));
   BUFX6TS FE_OCPUNCOC1070_FE_OFN377_offset_21_ (.Y(FE_OCPUNCON1070_FE_OFN377_offset_21_), 
	.A(FE_OFN377_offset_21_));
   BUFX16TS FE_OCPUNCOC1069_FE_OFN369_offset_23_ (.Y(FE_OCPUNCON1069_FE_OFN369_offset_23_), 
	.A(FE_OFN369_offset_23_));
   BUFX20TS FE_OCPUNCOC1068_offset_0_ (.Y(FE_OCPUNCON1068_offset_0_), 
	.A(offset[0]));
   BUFX20TS FE_OCPUNCOC1065_offset_2_ (.Y(FE_OCPUNCON1065_offset_2_), 
	.A(offset[2]));
   BUFX20TS FE_OCPUNCOC1060_offset_21_ (.Y(FE_OCPUNCON1060_offset_21_), 
	.A(offset[21]));
   CLKBUFX3TS FE_OCPUNCOC1058_filesize_3_ (.Y(FE_OCPUNCON1058_filesize_3_), 
	.A(filesize[3]));
   XNOR2X4TS FE_RC_417_0 (.Y(FE_OFN133_addr_calc_fft_read_addr_28_), 
	.B(\add_x_19_0/n4 ), 
	.A(\add_x_19_0/n50 ));
   XNOR2X4TS FE_RC_416_0 (.Y(FE_OFN135_addr_calc_fft_read_addr_30_), 
	.B(n1544), 
	.A(\add_x_19_0/n38 ));
   XNOR2X4TS FE_RC_415_0 (.Y(FE_OFN125_addr_calc_iir_write_addr_19_), 
	.B(\add_x_19_5/n13 ), 
	.A(\add_x_19_5/n99 ));
   XNOR2X4TS FE_RC_414_0 (.Y(FE_OFN123_addr_calc_iir_write_addr_21_), 
	.B(\add_x_19_5/n11 ), 
	.A(\add_x_19_5/n88 ));
   XNOR2X4TS FE_RC_413_0 (.Y(FE_OFN136_addr_calc_fft_read_addr_29_), 
	.B(n1451), 
	.A(FE_OCPN1730_add_x_19_0_n43));
   XNOR2X4TS FE_RC_412_0 (.Y(FE_OFN124_addr_calc_iir_write_addr_16_), 
	.B(\add_x_19_5/n16 ), 
	.A(\add_x_19_5/n112 ));
   XNOR2X4TS FE_RC_411_0 (.Y(FE_OFN128_addr_calc_iir_write_addr_10_), 
	.B(\add_x_19_5/n22 ), 
	.A(\add_x_19_5/n146 ));
   XNOR2X4TS FE_RC_410_0 (.Y(FE_OFN127_addr_calc_iir_write_addr_9_), 
	.B(\add_x_19_5/n23 ), 
	.A(\add_x_19_5/n153 ));
   OAI21X4TS FE_RC_408_0 (.Y(FE_OFN140_add_x_19_5_n115), 
	.B0(FE_RN_112_0), 
	.A1(\add_x_19_5/n116 ), 
	.A0(\add_x_19_5/n136 ));
   NAND2X8TS FE_RC_407_0 (.Y(FE_OFN139_add_x_19_0_n157), 
	.B(FE_RN_102_0), 
	.A(FE_RN_100_0));
   OR2X4TS FE_RC_390_0 (.Y(FE_RN_184_0), 
	.B(\add_x_19_0/n139 ), 
	.A(n1312));
   INVX2TS FE_RC_389_0 (.Y(FE_RN_183_0), 
	.A(\add_x_19_0/n139 ));
   CLKINVX1TS FE_RC_388_0 (.Y(FE_RN_182_0), 
	.A(n1312));
   OAI2BB1X2TS FE_RC_387_0 (.Y(FE_RN_181_0), 
	.B0(n1311), 
	.A1N(FE_RN_182_0), 
	.A0N(FE_RN_183_0));
   OAI21X2TS FE_RC_386_0 (.Y(\addr_calc/fft_read_addr[11] ), 
	.B0(FE_RN_181_0), 
	.A1(FE_RN_184_0), 
	.A0(n1311));
   NAND2X2TS FE_RC_380_0 (.Y(FE_RN_176_0), 
	.B(\add_x_19_2/n160 ), 
	.A(\add_x_19_2/n168 ));
   INVX2TS FE_RC_379_0 (.Y(FE_RN_175_0), 
	.A(\add_x_19_2/n169 ));
   INVX2TS FE_RC_378_0 (.Y(FE_RN_174_0), 
	.A(\add_x_19_2/n160 ));
   OA21X4TS FE_RC_377_0 (.Y(FE_RN_173_0), 
	.B0(\add_x_19_2/n163 ), 
	.A1(\add_x_19_2/n166 ), 
	.A0(\add_x_19_2/n162 ));
   OAI21X4TS FE_RC_371_0 (.Y(\add_x_19_5/n80 ), 
	.B0(\add_x_19_5/n82 ), 
	.A1(\add_x_19_5/n81 ), 
	.A0(\add_x_19_5/n83 ));
   OAI2BB1X2TS FE_RC_367_0 (.Y(\addr_calc/fir_read_addr[18] ), 
	.B0(FE_RN_135_0), 
	.A1N(\add_x_19_2/n102 ), 
	.A0N(FE_RN_136_0));
   INVX2TS FE_RC_366_0 (.Y(FE_RN_168_0), 
	.A(\add_x_19_4/n15 ));
   NAND2BX4TS FE_RC_365_0 (.Y(FE_RN_167_0), 
	.B(\add_x_19_4/n15 ), 
	.AN(\add_x_19_4/n107 ));
   OAI2BB1X4TS FE_RC_364_0 (.Y(\addr_calc/iir_read_addr[17] ), 
	.B0(FE_RN_167_0), 
	.A1N(\add_x_19_4/n107 ), 
	.A0N(FE_RN_168_0));
   XOR2X4TS FE_RC_363_0 (.Y(\addr_calc/fir_write_addr[22] ), 
	.B(n1391), 
	.A(\add_x_19_3/n83 ));
   XNOR2X4TS FE_RC_362_0 (.Y(\addr_calc/fft_read_addr[16] ), 
	.B(n1420), 
	.A(\add_x_19_0/n112 ));
   NAND2X2TS FE_RC_361_0 (.Y(FE_RN_166_0), 
	.B(n1605), 
	.A(\add_x_19_5/n60 ));
   NAND2X2TS FE_RC_360_0 (.Y(n1604), 
	.B(n1606), 
	.A(FE_RN_166_0));
   AOI21X4TS FE_RC_356_0 (.Y(\add_x_19_4/n83 ), 
	.B0(\add_x_19_4/n85 ), 
	.A1(\add_x_19_4/n84 ), 
	.A0(\add_x_19_4/n92 ));
   OAI21X2TS FE_RC_353_0 (.Y(\add_x_19_5/n130 ), 
	.B0(\add_x_19_5/n132 ), 
	.A1(\add_x_19_5/n131 ), 
	.A0(\add_x_19_5/n133 ));
   OAI21X4TS FE_RC_351_0 (.Y(\add_x_19_3/n146 ), 
	.B0(\add_x_19_3/n148 ), 
	.A1(\add_x_19_3/n147 ), 
	.A0(\add_x_19_3/n156 ));
   INVX2TS FE_RC_350_0 (.Y(FE_RN_165_0), 
	.A(\add_x_19_2/n44 ));
   NAND2BX4TS FE_RC_349_0 (.Y(FE_RN_164_0), 
	.B(FE_RN_165_0), 
	.AN(FE_OFN526_add_x_19_2_n113));
   NAND2X6TS FE_RC_348_0 (.Y(\add_x_19_2/n43 ), 
	.B(\add_x_19_2/n45 ), 
	.A(FE_RN_164_0));
   AOI21X4TS FE_RC_347_0 (.Y(\add_x_19_4/n125 ), 
	.B0(\add_x_19_4/n127 ), 
	.A1(\add_x_19_4/n126 ), 
	.A0(\add_x_19_4/n134 ));
   AOI21X4TS FE_RC_345_0 (.Y(\add_x_19_4/n136 ), 
	.B0(\add_x_19_4/n138 ), 
	.A1(\add_x_19_4/n137 ), 
	.A0(\add_x_19_4/n150 ));
   OAI21X2TS FE_RC_343_0 (.Y(\add_x_19_4/n150 ), 
	.B0(\add_x_19_4/n152 ), 
	.A1(\add_x_19_4/n151 ), 
	.A0(\add_x_19_4/n155 ));
   INVX2TS FE_RC_339_0 (.Y(FE_RN_163_0), 
	.A(\add_x_19_5/n180 ));
   OAI2BB1X4TS FE_RC_338_0 (.Y(n1818), 
	.B0(FE_RN_163_0), 
	.A1N(\add_x_19_5/n179 ), 
	.A0N(FE_OCPN1907_add_x_19_5_n187));
   INVX2TS FE_RC_336_0 (.Y(FE_RN_162_0), 
	.A(\add_x_19_5/n9 ));
   NAND2BX4TS FE_RC_335_0 (.Y(FE_RN_161_0), 
	.B(FE_RN_162_0), 
	.AN(\add_x_19_5/n80 ));
   INVX2TS FE_RC_330_0 (.Y(FE_RN_158_0), 
	.A(\add_x_19_5/n85 ));
   OAI2BB1X4TS FE_RC_329_0 (.Y(FE_RN_132_0), 
	.B0(FE_RN_158_0), 
	.A1N(\add_x_19_5/n92 ), 
	.A0N(\add_x_19_5/n84 ));
   INVX2TS FE_RC_328_0 (.Y(FE_RN_157_0), 
	.A(\add_x_19_2/n42 ));
   NAND2X2TS FE_RC_326_0 (.Y(FE_RN_156_0), 
	.B(\add_x_19_1/n46 ), 
	.A(\add_x_19_1/n72 ));
   OAI21X2TS FE_RC_325_0 (.Y(FE_RN_155_0), 
	.B0(\add_x_19_1/n49 ), 
	.A1(\add_x_19_1/n48 ), 
	.A0(\add_x_19_1/n52 ));
   AOI21X2TS FE_RC_324_0 (.Y(FE_RN_154_0), 
	.B0(FE_RN_155_0), 
	.A1(\add_x_19_1/n46 ), 
	.A0(\add_x_19_1/n73 ));
   OAI21X4TS FE_RC_323_0 (.Y(\add_x_19_1/n43 ), 
	.B0(FE_RN_154_0), 
	.A1(FE_RN_156_0), 
	.A0(FE_OFN523_add_x_19_1_n113));
   OAI21X1TS FE_RC_322_0 (.Y(FE_RN_153_0), 
	.B0(\add_x_19_1/n79 ), 
	.A1(\add_x_19_1/n82 ), 
	.A0(\add_x_19_1/n78 ));
   AOI21X2TS FE_RC_321_0 (.Y(FE_RN_152_0), 
	.B0(FE_RN_153_0), 
	.A1(\add_x_19_1/n85 ), 
	.A0(\add_x_19_1/n76 ));
   OR2X2TS FE_RC_315_0 (.Y(FE_RN_149_0), 
	.B(n2588), 
	.A(FE_OFN332_data_cntl_N63));
   OR3X8TS FE_RC_314_0 (.Y(n1701), 
	.C(FE_RN_149_0), 
	.B(n2793), 
	.A(n783));
   INVX2TS FE_RC_309_0 (.Y(FE_RN_146_0), 
	.A(n1949));
   INVX2TS FE_RC_308_0 (.Y(FE_RN_145_0), 
	.A(n1949));
   NAND2X4TS FE_RC_307_0 (.Y(FE_RN_144_0), 
	.B(FE_RN_145_0), 
	.A(n1730));
   OAI21X2TS FE_RC_306_0 (.Y(\DP_OP_158_296_6262/n1027 ), 
	.B0(FE_RN_144_0), 
	.A1(FE_RN_146_0), 
	.A0(n1730));
   XOR2X4TS FE_RC_305_0 (.Y(\addr_calc/iir_write_addr[22] ), 
	.B(n1323), 
	.A(\add_x_19_5/n83 ));
   CLKINVX1TS FE_RC_304_0 (.Y(FE_RN_143_0), 
	.A(n1434));
   NAND2BX2TS FE_RC_303_0 (.Y(FE_RN_142_0), 
	.B(n1434), 
	.AN(\add_x_19_0/n83 ));
   OAI2BB1X4TS FE_RC_302_0 (.Y(\addr_calc/fft_read_addr[22] ), 
	.B0(FE_RN_142_0), 
	.A1N(\add_x_19_0/n83 ), 
	.A0N(FE_RN_143_0));
   AOI21X4TS FE_RC_292_0 (.Y(\add_x_19_0/n60 ), 
	.B0(\add_x_19_0/n62 ), 
	.A1(\add_x_19_0/n61 ), 
	.A0(\add_x_19_0/n69 ));
   XOR2X4TS FE_RC_290_0 (.Y(\addr_calc/iir_read_addr[20] ), 
	.B(n1279), 
	.A(\add_x_19_4/n91 ));
   XOR2X4TS FE_RC_289_0 (.Y(\addr_calc/fir_write_addr[18] ), 
	.B(n1431), 
	.A(\add_x_19_3/n102 ));
   XOR2X4TS FE_RC_287_0 (.Y(\addr_calc/fir_read_addr[30] ), 
	.B(n1277), 
	.A(\add_x_19_2/n38 ));
   OAI2BB1X4TS FE_RC_286_0 (.Y(\add_x_19_3/n43 ), 
	.B0(n1299), 
	.A1N(FE_OCP_RBN1378_add_x_19_3_n113), 
	.A0N(n1470));
   CLKINVX1TS FE_RC_285_0 (.Y(FE_RN_136_0), 
	.A(n1432));
   NAND2BX2TS FE_RC_284_0 (.Y(FE_RN_135_0), 
	.B(n1432), 
	.AN(\add_x_19_2/n102 ));
   XNOR2X4TS FE_RC_281_0 (.Y(\addr_calc/fir_read_addr[16] ), 
	.B(n1416), 
	.A(\add_x_19_2/n112 ));
   AOI21X4TS FE_RC_278_0 (.Y(\add_x_19_5/n136 ), 
	.B0(\add_x_19_5/n138 ), 
	.A1(\add_x_19_5/n137 ), 
	.A0(\add_x_19_5/n150 ));
   OAI21X2TS FE_RC_277_0 (.Y(\add_x_19_5/n150 ), 
	.B0(\add_x_19_5/n152 ), 
	.A1(\add_x_19_5/n155 ), 
	.A0(\add_x_19_5/n151 ));
   INVX2TS FE_RC_276_0 (.Y(FE_RN_134_0), 
	.A(\add_x_19_3/n42 ));
   AOI21X4TS FE_RC_275_0 (.Y(\add_x_19_3/n38 ), 
	.B0(FE_RN_134_0), 
	.A1(n2631), 
	.A0(\add_x_19_3/n43 ));
   INVX8TS FE_RC_273_0 (.Y(\add_x_19_5/n83 ), 
	.A(FE_RN_132_0));
   INVX2TS FE_RC_267_0 (.Y(FE_RN_129_0), 
	.A(\add_x_19_0/n72 ));
   INVX2TS FE_RC_266_0 (.Y(FE_RN_128_0), 
	.A(\add_x_19_0/n73 ));
   OAI21X4TS FE_RC_265_0 (.Y(\add_x_19_0/n69 ), 
	.B0(FE_RN_128_0), 
	.A1(FE_RN_129_0), 
	.A0(FE_OFN528_add_x_19_0_n113));
   OAI21X2TS FE_RC_246_0 (.Y(FE_RN_113_0), 
	.B0(\add_x_19_5/n121 ), 
	.A1(\add_x_19_5/n120 ), 
	.A0(\add_x_19_5/n124 ));
   AOI21X4TS FE_RC_245_0 (.Y(FE_RN_112_0), 
	.B0(FE_RN_113_0), 
	.A1(\add_x_19_5/n127 ), 
	.A0(\add_x_19_5/n118 ));
   INVX3TS FE_RC_242_0 (.Y(FE_RN_110_0), 
	.A(\add_x_19_3/n178 ));
   NAND2X6TS FE_RC_240_0 (.Y(FE_RN_108_0), 
	.B(\add_x_19_3/n160 ), 
	.A(\add_x_19_3/n169 ));
   NAND2X4TS FE_RC_238_0 (.Y(FE_RN_107_0), 
	.B(\add_x_19_5/n160 ), 
	.A(\add_x_19_5/n168 ));
   OAI21X2TS FE_RC_233_0 (.Y(FE_RN_103_0), 
	.B0(\add_x_19_0/n163 ), 
	.A1(\add_x_19_0/n166 ), 
	.A0(\add_x_19_0/n162 ));
   AOI21X4TS FE_RC_232_0 (.Y(FE_RN_102_0), 
	.B0(FE_RN_103_0), 
	.A1(n1558), 
	.A0(\add_x_19_0/n169 ));
   INVX3TS FE_RC_231_0 (.Y(FE_RN_101_0), 
	.A(\add_x_19_0/n178 ));
   OAI21X2TS FE_RC_228_0 (.Y(FE_RN_99_0), 
	.B0(\add_x_19_0/n140 ), 
	.A1(\add_x_19_0/n145 ), 
	.A0(\add_x_19_0/n139 ));
   OAI21X1TS FE_RC_226_0 (.Y(FE_RN_98_0), 
	.B0(\add_x_19_2/n140 ), 
	.A1(\add_x_19_2/n145 ), 
	.A0(\add_x_19_2/n139 ));
   AOI21X4TS FE_RC_225_0 (.Y(\add_x_19_2/n136 ), 
	.B0(FE_RN_98_0), 
	.A1(\add_x_19_2/n137 ), 
	.A0(\add_x_19_2/n150 ));
   OAI21X2TS FE_RC_221_0 (.Y(\add_x_19_5/n88 ), 
	.B0(\add_x_19_5/n90 ), 
	.A1(\add_x_19_5/n89 ), 
	.A0(\add_x_19_5/n91 ));
   OAI21X4TS FE_RC_220_0 (.Y(\add_x_19_0/n99 ), 
	.B0(\add_x_19_0/n101 ), 
	.A1(\add_x_19_0/n102 ), 
	.A0(\add_x_19_0/n100 ));
   OAI21X4TS FE_RC_219_0 (.Y(\add_x_19_0/n88 ), 
	.B0(\add_x_19_0/n90 ), 
	.A1(\add_x_19_0/n89 ), 
	.A0(FE_OCP_RBN1383_add_x_19_0_n92));
   OAI21X2TS FE_RC_218_0 (.Y(n1300), 
	.B0(\add_x_19_3/n132 ), 
	.A1(\add_x_19_3/n131 ), 
	.A0(\add_x_19_3/n133 ));
   XOR2X4TS FE_RC_213_0 (.Y(\addr_calc/fft_read_addr[18] ), 
	.B(n1351), 
	.A(\add_x_19_0/n102 ));
   XOR2X4TS FE_RC_211_0 (.Y(\addr_calc/iir_write_addr[18] ), 
	.B(n1387), 
	.A(\add_x_19_5/n102 ));
   CLKINVX1TS FE_RC_210_0 (.Y(FE_RN_92_0), 
	.A(n1388));
   NAND2BX2TS FE_RC_209_0 (.Y(FE_RN_91_0), 
	.B(n1388), 
	.AN(\add_x_19_4/n102 ));
   OAI2BB1X4TS FE_RC_208_0 (.Y(\addr_calc/iir_read_addr[18] ), 
	.B0(FE_RN_91_0), 
	.A1N(\add_x_19_4/n102 ), 
	.A0N(FE_RN_92_0));
   XNOR2X4TS FE_RC_207_0 (.Y(\addr_calc/iir_write_addr[29] ), 
	.B(n1408), 
	.A(FE_OFN531_add_x_19_5_n43));
   XNOR2X4TS FE_RC_201_0 (.Y(\addr_calc/fft_write_addr[16] ), 
	.B(n1447), 
	.A(\add_x_19_1/n112 ));
   AOI21X4TS FE_RC_200_0 (.Y(\add_x_19_5/n60 ), 
	.B0(\add_x_19_5/n62 ), 
	.A1(\add_x_19_5/n61 ), 
	.A0(\add_x_19_5/n69 ));
   AOI21X4TS FE_RC_197_0 (.Y(\add_x_19_4/n159 ), 
	.B0(\add_x_19_4/n161 ), 
	.A1(\add_x_19_4/n160 ), 
	.A0(\add_x_19_4/n169 ));
   OR2X2TS FE_RC_194_0 (.Y(FE_RN_87_0), 
	.B(\add_x_19_4/n151 ), 
	.A(n1410));
   OR2X2TS FE_RC_193_0 (.Y(FE_RN_86_0), 
	.B(n1410), 
	.A(\add_x_19_4/n151 ));
   CLKINVX4TS FE_RC_191_0 (.Y(FE_RN_85_0), 
	.A(\add_x_19_5/n72 ));
   INVX2TS FE_RC_190_0 (.Y(FE_RN_84_0), 
	.A(\add_x_19_5/n73 ));
   OAI21X4TS FE_RC_189_0 (.Y(\add_x_19_5/n69 ), 
	.B0(FE_RN_84_0), 
	.A1(FE_RN_85_0), 
	.A0(\add_x_19_5/n113 ));
   OAI21X2TS FE_RC_164_0 (.Y(FE_RN_64_0), 
	.B0(\add_x_19_0/n98 ), 
	.A1(\add_x_19_0/n101 ), 
	.A0(\add_x_19_0/n97 ));
   OAI21X2TS FE_RC_157_0 (.Y(FE_RN_59_0), 
	.B0(\add_x_19_3/n98 ), 
	.A1(\add_x_19_3/n101 ), 
	.A0(\add_x_19_3/n97 ));
   AOI21X4TS FE_RC_156_0 (.Y(\add_x_19_3/n94 ), 
	.B0(FE_RN_59_0), 
	.A1(\add_x_19_3/n95 ), 
	.A0(\add_x_19_3/n104 ));
   NAND2X2TS FE_RC_152_0 (.Y(FE_RN_56_0), 
	.B(n2039), 
	.A(FE_OCPUNCON1576_n2812));
   NAND2X2TS FE_RC_151_0 (.Y(FE_RN_55_0), 
	.B(\addr_calc/iir_write_calc/counter/N49 ), 
	.A(FE_OCPUNCON1888_n2813));
   NAND2X2TS FE_RC_150_0 (.Y(n996), 
	.B(FE_RN_56_0), 
	.A(FE_RN_55_0));
   AOI21X4TS FE_RC_137_0 (.Y(n2812), 
	.B0(n1861), 
	.A1(FE_OFN315_data_from_iir), 
	.A0(\addr_calc/iir_write_calc/counter/N38 ));
   INVX2TS FE_RC_136_0 (.Y(FE_RN_46_0), 
	.A(\add_x_19_0/n11 ));
   NAND2BX2TS FE_RC_135_0 (.Y(FE_RN_45_0), 
	.B(FE_RN_46_0), 
	.AN(\add_x_19_0/n88 ));
   OAI2BB1X4TS FE_RC_134_0 (.Y(\addr_calc/fft_read_addr[21] ), 
	.B0(FE_RN_45_0), 
	.A1N(\add_x_19_0/n88 ), 
	.A0N(\add_x_19_0/n11 ));
   XOR2X4TS FE_RC_130_0 (.Y(\addr_calc/fir_write_addr[24] ), 
	.B(n1334), 
	.A(FE_OCPN1825_add_x_19_3_n68));
   XOR2X4TS FE_RC_129_0 (.Y(\DP_OP_159_297_3515/n51 ), 
	.B(\addr_calc/iir_read_calc/count[28] ), 
	.A(\DP_OP_159_297_3515/n1138 ));
   NOR2X1TS FE_RC_123_0 (.Y(FE_RN_41_0), 
	.B(\add_x_19_3/n151 ), 
	.A(n1283));
   NAND2BX2TS FE_RC_122_0 (.Y(FE_RN_40_0), 
	.B(FE_RN_41_0), 
	.AN(n1282));
   NAND2X4TS FE_RC_121_0 (.Y(\addr_calc/fir_write_addr[9] ), 
	.B(n1284), 
	.A(FE_RN_40_0));
   OAI2BB1X4TS FE_RC_120_0 (.Y(n1331), 
	.B0(\add_x_19_3/n111 ), 
	.A1N(FE_OCP_RBN1378_add_x_19_3_n113), 
	.A0N(\add_x_19_3/n207 ));
   XOR2X4TS FE_RC_119_0 (.Y(\addr_calc/iir_write_addr[14] ), 
	.B(n1360), 
	.A(\add_x_19_5/n125 ));
   OAI21X2TS FE_RC_118_0 (.Y(\add_x_19_3/n92 ), 
	.B0(\add_x_19_3/n94 ), 
	.A1(\add_x_19_3/n93 ), 
	.A0(\add_x_19_3/n113 ));
   INVX2TS FE_RC_117_0 (.Y(FE_RN_39_0), 
	.A(\add_x_19_3/n151 ));
   CLKINVX1TS FE_RC_116_0 (.Y(FE_RN_38_0), 
	.A(n1283));
   OAI2BB1X1TS FE_RC_115_0 (.Y(n1284), 
	.B0(n1282), 
	.A1N(FE_RN_38_0), 
	.A0N(FE_RN_39_0));
   OAI21X4TS FE_RC_113_0 (.Y(\add_x_19_3/n134 ), 
	.B0(FE_OCPN1908_add_x_19_3_n136), 
	.A1(\add_x_19_3/n135 ), 
	.A0(\add_x_19_3/n156 ));
   OAI21X2TS FE_RC_112_0 (.Y(\add_x_19_0/n146 ), 
	.B0(\add_x_19_0/n148 ), 
	.A1(\add_x_19_0/n147 ), 
	.A0(\add_x_19_0/n156 ));
   AOI21X4TS FE_RC_110_0 (.Y(\add_x_19_0/n117 ), 
	.B0(\add_x_19_0/n119 ), 
	.A1(\add_x_19_0/n118 ), 
	.A0(\add_x_19_0/n127 ));
   INVX8TS FE_RC_102_0 (.Y(\add_x_19_0/n112 ), 
	.A(FE_OCPN1728_FE_OFN528_add_x_19_0_n113));
   INVX2TS FE_RC_101_0 (.Y(FE_RN_35_0), 
	.A(\add_x_19_0/n207 ));
   NAND2BX4TS FE_RC_100_0 (.Y(FE_RN_34_0), 
	.B(FE_RN_35_0), 
	.AN(\add_x_19_0/n109 ));
   INVX2TS FE_RC_99_0 (.Y(FE_RN_33_0), 
	.A(\add_x_19_0/n109 ));
   NAND2X8TS FE_RC_98_0 (.Y(FE_RN_32_0), 
	.B(FE_RN_33_0), 
	.A(FE_OCPN1729_FE_OFN528_add_x_19_0_n113));
   NAND2X4TS FE_RC_97_0 (.Y(\add_x_19_0/n107 ), 
	.B(FE_RN_34_0), 
	.A(FE_RN_32_0));
   INVX2TS FE_RC_95_0 (.Y(FE_RN_31_0), 
	.A(\add_x_19_0/n127 ));
   OAI2BB1X4TS FE_RC_94_0 (.Y(FE_RN_30_0), 
	.B0(\add_x_19_0/n126 ), 
	.A1N(\add_x_19_0/n135 ), 
	.A0N(\add_x_19_0/n136 ));
   INVX2TS FE_RC_93_0 (.Y(FE_RN_29_0), 
	.A(\add_x_19_0/n127 ));
   NAND3X2TS FE_RC_92_0 (.Y(FE_RN_28_0), 
	.C(FE_RN_29_0), 
	.B(\add_x_19_0/n136 ), 
	.A(\add_x_19_0/n156 ));
   OAI2BB1X4TS FE_RC_91_0 (.Y(\add_x_19_0/n125 ), 
	.B0(FE_RN_28_0), 
	.A1N(FE_RN_30_0), 
	.A0N(FE_RN_31_0));
   CLKINVX12TS FE_RC_55_0 (.Y(n2441), 
	.A(FE_OCP_RBN1364_FE_OCP_DRV_N1167_offset_20_));
   INVX8TS FE_RC_54_0 (.Y(FE_OFN557_n2441), 
	.A(FE_OCP_RBN1364_FE_OCP_DRV_N1167_offset_20_));
   CLKINVX12TS FE_RC_53_0 (.Y(FE_OFN558_n2441), 
	.A(FE_OCP_RBN1366_FE_OCP_DRV_N1167_offset_20_));
   INVX2TS FE_RC_52_0 (.Y(FE_RN_7_0), 
	.A(n2048));
   AND2X8TS FE_RC_51_0 (.Y(\add_x_19_5/n89 ), 
	.B(FE_OCP_RBN1365_FE_OCP_DRV_N1167_offset_20_), 
	.A(FE_RN_7_0));
   BUFX20TS FE_RC_50_0 (.Y(FE_OFN411_offset_12_), 
	.A(FE_OFN410_offset_12_));
   BUFX20TS FE_RC_49_0 (.Y(FE_OFN413_offset_12_), 
	.A(FE_OFN410_offset_12_));
   CLKINVX4TS FE_RC_48_0 (.Y(\add_x_19_0/n131 ), 
	.A(FE_RN_5_0));
   INVX2TS FE_RC_47_0 (.Y(FE_RN_6_0), 
	.A(n2046));
   NAND2BX4TS FE_RC_46_0 (.Y(FE_RN_5_0), 
	.B(FE_RN_6_0), 
	.AN(FE_OFN410_offset_12_));
   NOR2BX4TS FE_RC_45_0 (.Y(\add_x_19_0/n126 ), 
	.B(\add_x_19_0/n128 ), 
	.AN(FE_RN_5_0));
   BUFX20TS FE_RC_39_0 (.Y(FE_OFN418_offset_10_), 
	.A(offset[10]));
   BUFX20TS FE_RC_38_0 (.Y(FE_OCPUNCON653_FE_OFN418_offset_10_), 
	.A(offset[10]));
   BUFX20TS FE_RC_37_0 (.Y(FE_OCPUNCON657_FE_OFN418_offset_10_), 
	.A(offset[10]));
   NOR2X1TS FE_RC_36_0 (.Y(\add_x_19_0/n144 ), 
	.B(offset[10]), 
	.A(\addr_calc/fft_read_calc/count[10] ));
   BUFX20TS FE_RC_34_0 (.Y(FE_OFN435_offset_6_), 
	.A(offset[6]));
   BUFX20TS FE_RC_33_0 (.Y(FE_OCPUNCON726_FE_OFN435_offset_6_), 
	.A(offset[6]));
   CLKINVX4TS FE_RC_32_0 (.Y(\add_x_19_3/n165 ), 
	.A(FE_RN_1_0));
   INVX2TS FE_RC_31_0 (.Y(FE_RN_2_0), 
	.A(FE_OFN253_addr_calc_fir_write_calc_count_6_));
   NAND2BX4TS FE_RC_30_0 (.Y(FE_RN_1_0), 
	.B(FE_RN_2_0), 
	.AN(offset[6]));
   NOR2BX4TS FE_RC_29_0 (.Y(\add_x_19_3/n160 ), 
	.B(\add_x_19_3/n162 ), 
	.AN(FE_RN_1_0));
   BUFX20TS FE_RC_27_0 (.Y(FE_OFN461_offset_0_), 
	.A(offset[0]));
   NAND2X1TS FE_RC_26_0 (.Y(\add_x_19_0/n191 ), 
	.B(n2058), 
	.A(offset[0]));
   NAND2X8TS FE_RC_25_0 (.Y(FE_RN_0_0), 
	.B(offset[0]), 
	.A(n2058));
   OAI21X4TS FE_RC_24_0 (.Y(\add_x_19_0/n187 ), 
	.B0(\add_x_19_0/n189 ), 
	.A1(\add_x_19_0/n188 ), 
	.A0(FE_RN_0_0));
   BUFX20TS FE_RC_23_0 (.Y(FE_OCPUNCON654_FE_OFN422_offset_9_), 
	.A(FE_OFN422_offset_9_));
   BUFX20TS FE_RC_22_0 (.Y(FE_OCPUNCON658_FE_OFN422_offset_9_), 
	.A(FE_OFN422_offset_9_));
   NOR2X8TS FE_RC_19_0 (.Y(\add_x_19_0/n188 ), 
	.B(FE_OCPUNCON1750_offset_1_), 
	.A(\addr_calc/fft_read_calc/count[1] ));
   NOR2X8TS FE_RC_12_0 (.Y(\add_x_19_0/n181 ), 
	.B(\addr_calc/fft_read_calc/count[3] ), 
	.A(FE_OCPN1188_offset_3_));
   BUFX20TS FE_RC_10_0 (.Y(FE_OFN452_offset_2_), 
	.A(FE_OCPN1944_offset_2_));
   NOR2X8TS FE_RC_9_0 (.Y(\add_x_19_0/n184 ), 
	.B(FE_OCPN1945_offset_2_), 
	.A(\addr_calc/fft_read_calc/count[2] ));
   BUFX20TS FE_OCPUNCOC656_FE_OFN414_offset_11_ (.Y(FE_OCPUNCON656_FE_OFN414_offset_11_), 
	.A(FE_OCPUNCON652_FE_OFN414_offset_11_));
   BUFX20TS FE_OCPUNCOC652_FE_OFN414_offset_11_ (.Y(FE_OCPUNCON652_FE_OFN414_offset_11_), 
	.A(FE_OCPUNCON1873_offset_11_));
   BUFX3TS FE_OFC615_filesize_0_ (.Y(FE_OFN615_filesize_0_), 
	.A(FE_OCP_DRV_N1336_filesize_0_));
   CLKBUFX2TS FE_OFC612_filesize_4_ (.Y(FE_OFN612_filesize_4_), 
	.A(filesize[4]));
   CLKBUFX2TS FE_OFC611_filesize_5_ (.Y(FE_OFN611_filesize_5_), 
	.A(filesize[5]));
   CLKBUFX2TS FE_OFC610_filesize_6_ (.Y(FE_OFN610_filesize_6_), 
	.A(filesize[6]));
   CLKBUFX2TS FE_OFC609_filesize_7_ (.Y(FE_OFN609_filesize_7_), 
	.A(filesize[7]));
   BUFX3TS FE_OFC608_filesize_8_ (.Y(FE_OFN608_filesize_8_), 
	.A(FE_OCP_DRV_N1968_filesize_8_));
   CLKBUFX2TS FE_OFC607_filesize_9_ (.Y(FE_OFN607_filesize_9_), 
	.A(filesize[9]));
   CLKBUFX2TS FE_OFC605_filesize_11_ (.Y(FE_OFN605_filesize_11_), 
	.A(filesize[11]));
   CLKBUFX2TS FE_OFC604_filesize_12_ (.Y(FE_OFN604_filesize_12_), 
	.A(filesize[12]));
   CLKBUFX2TS FE_OFC603_filesize_13_ (.Y(FE_OFN603_filesize_13_), 
	.A(filesize[13]));
   BUFX3TS FE_OFC602_filesize_14_ (.Y(FE_OFN602_filesize_14_), 
	.A(FE_OCP_DRV_N1099_filesize_14_));
   CLKBUFX2TS FE_OFC600_filesize_17_ (.Y(FE_OFN600_filesize_17_), 
	.A(filesize[17]));
   BUFX3TS FE_OFC599_filesize_18_ (.Y(FE_OFN599_filesize_18_), 
	.A(FE_OCP_DRV_N1872_filesize_18_));
   BUFX3TS FE_OFC598_filesize_19_ (.Y(FE_OFN598_filesize_19_), 
	.A(FE_OCP_DRV_N1824_filesize_19_));
   BUFX3TS FE_OFC597_filesize_20_ (.Y(FE_OFN597_filesize_20_), 
	.A(FE_OCP_DRV_N1818_filesize_20_));
   CLKBUFX2TS FE_OFC596_filesize_21_ (.Y(FE_OFN596_filesize_21_), 
	.A(filesize[21]));
   CLKBUFX2TS FE_OFC595_filesize_24_ (.Y(FE_OFN595_filesize_24_), 
	.A(filesize[24]));
   CLKBUFX2TS FE_OFC594_filesize_26_ (.Y(FE_OFN594_filesize_26_), 
	.A(filesize[26]));
   CLKBUFX2TS FE_OFC593_filesize_27_ (.Y(FE_OFN593_filesize_27_), 
	.A(filesize[27]));
   CLKBUFX2TS FE_OFC592_filesize_28_ (.Y(FE_OFN592_filesize_28_), 
	.A(filesize[28]));
   BUFX3TS FE_OFC591_filesize_29_ (.Y(FE_OFN591_filesize_29_), 
	.A(FE_OCP_DRV_N1894_filesize_29_));
   CLKBUFX2TS FE_OFC567_n2070 (.Y(FE_OFN567_n2070), 
	.A(n2070));
   CLKBUFX2TS FE_OFC566_n2066 (.Y(FE_OFN566_n2066), 
	.A(FE_OFN565_n2066));
   CLKBUFX2TS FE_OFC565_n2066 (.Y(FE_OFN565_n2066), 
	.A(FE_OFN564_n2066));
   CLKBUFX2TS FE_OFC564_n2066 (.Y(FE_OFN564_n2066), 
	.A(n2066));
   CLKBUFX2TS FE_OFC563_n2060 (.Y(FE_OFN563_n2060), 
	.A(n2060));
   CLKBUFX2TS FE_OFC562_n2060 (.Y(FE_OFN562_n2060), 
	.A(n2060));
   CLKBUFX2TS FE_OFC561_n2587 (.Y(FE_OFN561_n2587), 
	.A(n2587));
   CLKBUFX2TS FE_OFC560_n2587 (.Y(FE_OFN560_n2587), 
	.A(n2587));
   CLKBUFX2TS FE_OFC559_offset_30_ (.Y(FE_OFN559_offset_30_), 
	.A(FE_OFN343_offset_30_));
   BUFX3TS FE_OFC553_n1789 (.Y(FE_OFN553_n1789), 
	.A(n1789));
   BUFX3TS FE_OFC552_n1751 (.Y(FE_OFN552_n1751), 
	.A(n1751));
   CLKBUFX2TS FE_OFC551_n1751 (.Y(FE_OFN551_n1751), 
	.A(FE_OFN1_n1751));
   CLKBUFX2TS FE_OFC550_n1750 (.Y(FE_OFN550_n1750), 
	.A(FE_OFN6_n1750));
   CLKBUFX2TS FE_OFC549_n1763 (.Y(FE_OFN549_n1763), 
	.A(n1763));
   CLKBUFX2TS FE_OFC548_n1763 (.Y(FE_OFN548_n1763), 
	.A(n1763));
   CLKBUFX3TS FE_OFC547_n2803 (.Y(FE_OFN547_n2803), 
	.A(n2803));
   BUFX8TS FE_OFC545_addr_calc_iir_write_addr_11_ (.Y(FE_OFN545_addr_calc_iir_write_addr_11_), 
	.A(\addr_calc/iir_write_addr[11] ));
   BUFX6TS FE_OFC544_addr_calc_fft_read_addr_11_ (.Y(FE_OFN544_addr_calc_fft_read_addr_11_), 
	.A(\addr_calc/fft_read_addr[11] ));
   BUFX6TS FE_OFC543_addr_calc_fir_write_addr_17_ (.Y(FE_OFN543_addr_calc_fir_write_addr_17_), 
	.A(\addr_calc/fir_write_addr[17] ));
   BUFX3TS FE_OFC540_DP_OP_158_296_6262_n765 (.Y(FE_OFN540_DP_OP_158_296_6262_n765), 
	.A(\DP_OP_158_296_6262/n765 ));
   BUFX4TS FE_OFC539_DP_OP_158_296_6262_n318 (.Y(FE_OFN539_DP_OP_158_296_6262_n318), 
	.A(\DP_OP_158_296_6262/n318 ));
   BUFX8TS FE_OFC538_DP_OP_158_296_6262_n1659 (.Y(FE_OFN538_DP_OP_158_296_6262_n1659), 
	.A(\DP_OP_158_296_6262/n1659 ));
   BUFX12TS FE_OFC537_DP_OP_159_297_3515_n301 (.Y(FE_OFN537_DP_OP_159_297_3515_n301), 
	.A(\DP_OP_159_297_3515/n301 ));
   BUFX8TS FE_OFC536_addr_calc_iir_read_addr_7_ (.Y(FE_OFN536_addr_calc_iir_read_addr_7_), 
	.A(\addr_calc/iir_read_addr[7] ));
   BUFX3TS FE_OFC535_DP_OP_159_297_3515_n726 (.Y(FE_OFN535_DP_OP_159_297_3515_n726), 
	.A(\DP_OP_159_297_3515/n726 ));
   BUFX6TS FE_OFC534_addr_calc_iir_write_addr_7_ (.Y(FE_OFN534_addr_calc_iir_write_addr_7_), 
	.A(\addr_calc/iir_write_addr[7] ));
   BUFX4TS FE_OFC533_addr_calc_fir_write_addr_7_ (.Y(FE_OFN533_addr_calc_fir_write_addr_7_), 
	.A(\addr_calc/fir_write_addr[7] ));
   BUFX6TS FE_OFC532_addr_calc_fft_read_addr_7_ (.Y(FE_OFN532_addr_calc_fft_read_addr_7_), 
	.A(\addr_calc/fft_read_addr[7] ));
   BUFX6TS FE_OFC531_add_x_19_5_n43 (.Y(FE_OFN531_add_x_19_5_n43), 
	.A(\add_x_19_5/n43 ));
   BUFX12TS FE_OFC529_DP_OP_158_296_6262_n838 (.Y(FE_OFN529_DP_OP_158_296_6262_n838), 
	.A(\DP_OP_158_296_6262/n838 ));
   BUFX16TS FE_OFC528_add_x_19_0_n113 (.Y(FE_OFN528_add_x_19_0_n113), 
	.A(\add_x_19_0/n113 ));
   BUFX16TS FE_OFC527_add_x_19_4_n113 (.Y(FE_OFN527_add_x_19_4_n113), 
	.A(\add_x_19_4/n113 ));
   BUFX16TS FE_OFC526_add_x_19_2_n113 (.Y(FE_OFN526_add_x_19_2_n113), 
	.A(\add_x_19_2/n113 ));
   BUFX4TS FE_OFC524_n1659 (.Y(FE_OFN524_n1659), 
	.A(n1659));
   BUFX16TS FE_OFC523_add_x_19_1_n113 (.Y(FE_OFN523_add_x_19_1_n113), 
	.A(\add_x_19_1/n113 ));
   BUFX8TS FE_OFC522_add_x_19_5_n114 (.Y(FE_OFN522_add_x_19_5_n114), 
	.A(\add_x_19_5/n114 ));
   BUFX12TS FE_OFC521_n1592 (.Y(FE_OFN521_n1592), 
	.A(n1592));
   BUFX20TS FE_OFC520_add_x_19_1_n157 (.Y(FE_OFN520_add_x_19_1_n157), 
	.A(\add_x_19_1/n157 ));
   BUFX12TS FE_OFC519_DP_OP_159_297_3515_n1039 (.Y(FE_OFN519_DP_OP_159_297_3515_n1039), 
	.A(\DP_OP_159_297_3515/n1039 ));
   BUFX3TS FE_OFC518_n2372 (.Y(FE_OFN518_n2372), 
	.A(n2372));
   CLKBUFX3TS FE_OFC517_addr_calc_fft_read_calc_count_0_ (.Y(FE_OFN517_addr_calc_fft_read_calc_count_0_), 
	.A(\addr_calc/fft_read_calc/count[0] ));
   CLKBUFX2TS FE_OFC516_from_iir_full (.Y(FE_OFN516_from_iir_full), 
	.A(from_iir_full));
   CLKBUFX2TS FE_OFC515_from_iir_empty (.Y(FE_OFN515_from_iir_empty), 
	.A(from_iir_empty));
   CLKBUFX2TS FE_OFC514_to_iir_full (.Y(FE_OFN514_to_iir_full), 
	.A(to_iir_full));
   CLKBUFX2TS FE_OFC513_to_iir_empty (.Y(FE_OFN513_to_iir_empty), 
	.A(to_iir_empty));
   CLKBUFX2TS FE_OFC512_from_fir_full (.Y(FE_OFN512_from_fir_full), 
	.A(from_fir_full));
   CLKBUFX2TS FE_OFC511_from_fir_empty (.Y(FE_OFN511_from_fir_empty), 
	.A(from_fir_empty));
   CLKBUFX2TS FE_OFC510_to_fir_full (.Y(FE_OFN510_to_fir_full), 
	.A(to_fir_full));
   CLKBUFX2TS FE_OFC509_to_fir_empty (.Y(FE_OFN509_to_fir_empty), 
	.A(to_fir_empty));
   CLKBUFX2TS FE_OFC508_from_fft_full (.Y(FE_OFN508_from_fft_full), 
	.A(from_fft_full));
   CLKBUFX2TS FE_OFC507_from_fft_empty (.Y(FE_OFN507_from_fft_empty), 
	.A(from_fft_empty));
   CLKBUFX2TS FE_OFC506_to_fft_full (.Y(FE_OFN506_to_fft_full), 
	.A(to_fft_full));
   CLKBUFX2TS FE_OFC505_to_fft_empty (.Y(FE_OFN505_to_fft_empty), 
	.A(to_fft_empty));
   CLKBUFX2TS FE_OFC504_iir_data_in_9_ (.Y(FE_OFN504_iir_data_in_9_), 
	.A(iir_data_in[9]));
   CLKBUFX2TS FE_OFC503_fft_data_in_9_ (.Y(FE_OFN503_fft_data_in_9_), 
	.A(fft_data_in[9]));
   BUFX20TS FE_OFC502_filesize_0_ (.Y(FE_OFN502_filesize_0_), 
	.A(FE_OFN615_filesize_0_));
   BUFX20TS FE_OFC501_filesize_1_ (.Y(FE_OFN501_filesize_1_), 
	.A(FE_OFN500_filesize_1_));
   BUFX20TS FE_OFC500_filesize_1_ (.Y(FE_OFN500_filesize_1_), 
	.A(FE_OFN614_filesize_1_));
   BUFX20TS FE_OFC499_filesize_2_ (.Y(FE_OFN499_filesize_2_), 
	.A(FE_OFN613_filesize_2_));
   BUFX8TS FE_OFC498_filesize_3_ (.Y(FE_OFN498_filesize_3_), 
	.A(FE_OCPUNCON1058_filesize_3_));
   CLKBUFX12TS FE_OFC496_filesize_4_ (.Y(FE_OFN496_filesize_4_), 
	.A(FE_OFN612_filesize_4_));
   BUFX20TS FE_OFC495_filesize_5_ (.Y(FE_OFN495_filesize_5_), 
	.A(FE_OFN611_filesize_5_));
   BUFX20TS FE_OFC494_filesize_6_ (.Y(FE_OFN494_filesize_6_), 
	.A(FE_OFN610_filesize_6_));
   BUFX20TS FE_OFC493_filesize_7_ (.Y(FE_OFN493_filesize_7_), 
	.A(FE_OFN609_filesize_7_));
   BUFX20TS FE_OFC492_filesize_8_ (.Y(FE_OFN492_filesize_8_), 
	.A(FE_OFN608_filesize_8_));
   BUFX16TS FE_OFC491_filesize_9_ (.Y(FE_OFN491_filesize_9_), 
	.A(FE_OFN607_filesize_9_));
   BUFX16TS FE_OFC490_filesize_10_ (.Y(FE_OFN490_filesize_10_), 
	.A(FE_OCPUNCON1562_filesize_10_));
   BUFX20TS FE_OFC489_filesize_11_ (.Y(FE_OFN489_filesize_11_), 
	.A(FE_OFN605_filesize_11_));
   BUFX20TS FE_OFC488_filesize_12_ (.Y(FE_OFN488_filesize_12_), 
	.A(FE_OFN604_filesize_12_));
   BUFX20TS FE_OFC487_filesize_13_ (.Y(FE_OFN487_filesize_13_), 
	.A(FE_OFN603_filesize_13_));
   BUFX20TS FE_OFC486_filesize_14_ (.Y(FE_OFN486_filesize_14_), 
	.A(FE_OFN485_filesize_14_));
   BUFX20TS FE_OFC485_filesize_14_ (.Y(FE_OFN485_filesize_14_), 
	.A(FE_OFN602_filesize_14_));
   BUFX8TS FE_OFC484_filesize_15_ (.Y(FE_OFN484_filesize_15_), 
	.A(FE_OFN483_filesize_15_));
   CLKBUFX3TS FE_OFC483_filesize_15_ (.Y(FE_OFN483_filesize_15_), 
	.A(filesize[15]));
   BUFX3TS FE_OFC482_filesize_16_ (.Y(FE_OFN482_filesize_16_), 
	.A(FE_OFN481_filesize_16_));
   BUFX20TS FE_OFC480_filesize_17_ (.Y(FE_OFN480_filesize_17_), 
	.A(FE_OFN600_filesize_17_));
   BUFX20TS FE_OFC479_filesize_18_ (.Y(FE_OFN479_filesize_18_), 
	.A(FE_OFN599_filesize_18_));
   BUFX20TS FE_OFC478_filesize_19_ (.Y(FE_OFN478_filesize_19_), 
	.A(FE_OFN598_filesize_19_));
   BUFX16TS FE_OFC477_filesize_20_ (.Y(FE_OFN477_filesize_20_), 
	.A(FE_OFN597_filesize_20_));
   CLKBUFX12TS FE_OFC476_filesize_21_ (.Y(FE_OFN476_filesize_21_), 
	.A(FE_OFN596_filesize_21_));
   BUFX8TS FE_OFC475_filesize_22_ (.Y(FE_OFN475_filesize_22_), 
	.A(FE_OFN474_filesize_22_));
   CLKBUFX3TS FE_OFC474_filesize_22_ (.Y(FE_OFN474_filesize_22_), 
	.A(filesize[22]));
   BUFX8TS FE_OFC473_filesize_23_ (.Y(FE_OFN473_filesize_23_), 
	.A(FE_OFN472_filesize_23_));
   CLKBUFX3TS FE_OFC472_filesize_23_ (.Y(FE_OFN472_filesize_23_), 
	.A(filesize[23]));
   BUFX20TS FE_OFC471_filesize_24_ (.Y(FE_OFN471_filesize_24_), 
	.A(FE_OFN595_filesize_24_));
   BUFX8TS FE_OFC470_filesize_25_ (.Y(FE_OFN470_filesize_25_), 
	.A(FE_OFN469_filesize_25_));
   CLKBUFX3TS FE_OFC469_filesize_25_ (.Y(FE_OFN469_filesize_25_), 
	.A(filesize[25]));
   BUFX20TS FE_OFC468_filesize_26_ (.Y(FE_OFN468_filesize_26_), 
	.A(FE_OFN594_filesize_26_));
   BUFX20TS FE_OFC467_filesize_27_ (.Y(FE_OFN467_filesize_27_), 
	.A(FE_OFN593_filesize_27_));
   BUFX20TS FE_OFC466_filesize_28_ (.Y(FE_OFN466_filesize_28_), 
	.A(FE_OFN592_filesize_28_));
   BUFX3TS FE_OFC465_filesize_29_ (.Y(FE_OFN465_filesize_29_), 
	.A(FE_OFN464_filesize_29_));
   BUFX20TS FE_OFC464_filesize_29_ (.Y(FE_OFN464_filesize_29_), 
	.A(FE_OFN591_filesize_29_));
   CLKBUFX3TS FE_OFC463_filesize_30_ (.Y(FE_OFN463_filesize_30_), 
	.A(filesize[30]));
   CLKBUFX3TS FE_OFC462_filesize_31_ (.Y(FE_OFN462_filesize_31_), 
	.A(filesize[31]));
   BUFX16TS FE_OFC459_offset_0_ (.Y(FE_OFN459_offset_0_), 
	.A(FE_OCPUNCON1068_offset_0_));
   BUFX20TS FE_OFC451_offset_2_ (.Y(FE_OFN451_offset_2_), 
	.A(FE_OCPUNCON1065_offset_2_));
   BUFX16TS FE_OFC447_offset_3_ (.Y(FE_OFN447_offset_3_), 
	.A(FE_OCPUNCON1066_offset_3_));
   BUFX8TS FE_OFC444_offset_4_ (.Y(FE_OFN444_offset_4_), 
	.A(FE_OCPUNCON1875_offset_4_));
   BUFX8TS FE_OFC443_offset_4_ (.Y(FE_OFN443_offset_4_), 
	.A(FE_OCPUNCON1875_offset_4_));
   BUFX16TS FE_OFC429_offset_8_ (.Y(FE_OFN429_offset_8_), 
	.A(FE_OFN427_offset_8_));
   BUFX16TS FE_OFC428_offset_8_ (.Y(FE_OFN428_offset_8_), 
	.A(FE_OFN426_offset_8_));
   BUFX20TS FE_OFC427_offset_8_ (.Y(FE_OFN427_offset_8_), 
	.A(FE_OFN426_offset_8_));
   BUFX20TS FE_OFC421_offset_10_ (.Y(FE_OFN421_offset_10_), 
	.A(FE_OFN418_offset_10_));
   CLKBUFX12TS FE_OFC417_offset_11_ (.Y(FE_OFN417_offset_11_), 
	.A(FE_OCPUNCON1873_offset_11_));
   CLKBUFX12TS FE_OFC408_offset_13_ (.Y(FE_OFN408_offset_13_), 
	.A(FE_OCPUNCON1941_offset_13_));
   BUFX16TS FE_OFC407_offset_13_ (.Y(FE_OFN407_offset_13_), 
	.A(FE_OCPUNCON1941_offset_13_));
   BUFX20TS FE_OFC400_offset_15_ (.Y(FE_OFN400_offset_15_), 
	.A(FE_OCPUNCON1940_offset_15_));
   BUFX16TS FE_OFC397_offset_16_ (.Y(FE_OFN397_offset_16_), 
	.A(FE_OFN395_offset_16_));
   BUFX20TS FE_OFC396_offset_16_ (.Y(FE_OFN396_offset_16_), 
	.A(FE_OFN394_offset_16_));
   BUFX16TS FE_OFC395_offset_16_ (.Y(FE_OFN395_offset_16_), 
	.A(FE_OFN394_offset_16_));
   BUFX20TS FE_OFC394_offset_16_ (.Y(FE_OFN394_offset_16_), 
	.A(FE_OFN580_offset_16_));
   BUFX16TS FE_OFC393_offset_17_ (.Y(FE_OFN393_offset_17_), 
	.A(FE_OFN391_offset_17_));
   BUFX8TS FE_OFC392_offset_17_ (.Y(FE_OFN392_offset_17_), 
	.A(FE_OFN390_offset_17_));
   BUFX16TS FE_OFC391_offset_17_ (.Y(FE_OFN391_offset_17_), 
	.A(FE_OFN390_offset_17_));
   CLKBUFX12TS FE_OFC389_offset_18_ (.Y(FE_OFN389_offset_18_), 
	.A(FE_OFN386_offset_18_));
   BUFX20TS FE_OFC384_offset_19_ (.Y(FE_OFN384_offset_19_), 
	.A(FE_OFN382_offset_19_));
   BUFX20TS FE_OFC382_offset_19_ (.Y(FE_OFN382_offset_19_), 
	.A(FE_OCPUNCON1062_offset_19_));
   BUFX20TS FE_OFC380_offset_21_ (.Y(FE_OFN380_offset_21_), 
	.A(FE_OFN377_offset_21_));
   BUFX20TS FE_OFC377_offset_21_ (.Y(FE_OFN377_offset_21_), 
	.A(FE_OCPUNCON1060_offset_21_));
   CLKBUFX12TS FE_OFC375_offset_22_ (.Y(FE_OFN375_offset_22_), 
	.A(FE_OCPUNCON1876_offset_22_));
   BUFX20TS FE_OFC374_offset_22_ (.Y(FE_OFN374_offset_22_), 
	.A(FE_OCPUNCON1876_offset_22_));
   BUFX8TS FE_OFC372_offset_23_ (.Y(FE_OFN372_offset_23_), 
	.A(FE_OCPUNCON1069_FE_OFN369_offset_23_));
   BUFX16TS FE_OFC371_offset_23_ (.Y(FE_OFN371_offset_23_), 
	.A(FE_OFN369_offset_23_));
   BUFX12TS FE_OFC368_offset_24_ (.Y(FE_OFN368_offset_24_), 
	.A(FE_OFN366_offset_24_));
   BUFX8TS FE_OFC367_offset_24_ (.Y(FE_OFN367_offset_24_), 
	.A(FE_OFN365_offset_24_));
   BUFX3TS FE_OFC366_offset_24_ (.Y(FE_OFN366_offset_24_), 
	.A(FE_OFN365_offset_24_));
   CLKBUFX12TS FE_OFC364_offset_25_ (.Y(FE_OFN364_offset_25_), 
	.A(FE_OFN361_offset_25_));
   BUFX8TS FE_OFC363_offset_25_ (.Y(FE_OFN363_offset_25_), 
	.A(FE_OCPUNCON1318_FE_OFN361_offset_25_));
   BUFX16TS FE_OFC360_offset_26_ (.Y(FE_OFN360_offset_26_), 
	.A(FE_OFN358_offset_26_));
   BUFX16TS FE_OFC359_offset_26_ (.Y(FE_OFN359_offset_26_), 
	.A(FE_OFN357_offset_26_));
   BUFX16TS FE_OFC358_offset_26_ (.Y(FE_OFN358_offset_26_), 
	.A(FE_OFN357_offset_26_));
   BUFX8TS FE_OFC356_offset_27_ (.Y(FE_OFN356_offset_27_), 
	.A(FE_OFN354_offset_27_));
   CLKBUFX12TS FE_OFC355_offset_27_ (.Y(FE_OFN355_offset_27_), 
	.A(FE_OFN353_offset_27_));
   BUFX3TS FE_OFC354_offset_27_ (.Y(FE_OFN354_offset_27_), 
	.A(FE_OFN353_offset_27_));
   BUFX8TS FE_OFC352_offset_28_ (.Y(FE_OFN352_offset_28_), 
	.A(FE_OFN350_offset_28_));
   CLKBUFX3TS FE_OFC351_offset_28_ (.Y(FE_OFN351_offset_28_), 
	.A(FE_OFN349_offset_28_));
   BUFX3TS FE_OFC350_offset_28_ (.Y(FE_OFN350_offset_28_), 
	.A(FE_OFN349_offset_28_));
   BUFX20TS FE_OFC349_offset_28_ (.Y(FE_OFN349_offset_28_), 
	.A(FE_OFN568_offset_28_));
   BUFX3TS FE_OFC348_offset_29_ (.Y(FE_OFN348_offset_29_), 
	.A(FE_OFN346_offset_29_));
   CLKBUFX2TS FE_OFC347_offset_29_ (.Y(FE_OFN347_offset_29_), 
	.A(FE_OFN345_offset_29_));
   CLKBUFX2TS FE_OFC346_offset_29_ (.Y(FE_OFN346_offset_29_), 
	.A(FE_OFN345_offset_29_));
   CLKBUFX3TS FE_OFC345_offset_29_ (.Y(FE_OFN345_offset_29_), 
	.A(offset[29]));
   CLKBUFX2TS FE_OFC344_offset_30_ (.Y(FE_OFN344_offset_30_), 
	.A(FE_OFN343_offset_30_));
   BUFX3TS FE_OFC343_offset_30_ (.Y(FE_OFN343_offset_30_), 
	.A(FE_OFN341_offset_30_));
   BUFX3TS FE_OFC341_offset_30_ (.Y(FE_OFN341_offset_30_), 
	.A(offset[30]));
   CLKBUFX2TS FE_OFC340_offset_31_ (.Y(FE_OFN340_offset_31_), 
	.A(FE_OFN338_offset_31_));
   CLKBUFX2TS FE_OFC339_offset_31_ (.Y(FE_OFN339_offset_31_), 
	.A(FE_OFN337_offset_31_));
   CLKBUFX2TS FE_OFC338_offset_31_ (.Y(FE_OFN338_offset_31_), 
	.A(FE_OFN337_offset_31_));
   CLKBUFX3TS FE_OFC337_offset_31_ (.Y(FE_OFN337_offset_31_), 
	.A(offset[31]));
   CLKBUFX2TS FE_OFC336_instruction_0_ (.Y(FE_OFN336_instruction_0_), 
	.A(instruction[0]));
   CLKBUFX2TS FE_OFC335_instruction_2_ (.Y(FE_OFN335_instruction_2_), 
	.A(instruction[2]));
   CLKBUFX2TS FE_OFC334_data_to_fft (.Y(FE_OFN334_data_to_fft), 
	.A(FE_OFN333_data_to_fft));
   CLKBUFX3TS FE_OFC333_data_to_fft (.Y(FE_OFN333_data_to_fft), 
	.A(data_to_fft));
   CLKBUFX3TS FE_OFC332_data_cntl_N63 (.Y(FE_OFN332_data_cntl_N63), 
	.A(\data_cntl/N63 ));
   CLKBUFX2TS FE_OFC331_data_to_fir (.Y(FE_OFN331_data_to_fir), 
	.A(FE_OFN330_data_to_fir));
   CLKBUFX2TS FE_OFC330_data_to_fir (.Y(FE_OFN330_data_to_fir), 
	.A(data_to_fir));
   CLKBUFX2TS FE_OFC329_data_cntl_N99 (.Y(FE_OFN329_data_cntl_N99), 
	.A(\data_cntl/N99 ));
   CLKBUFX2TS FE_OFC328_data_to_iir (.Y(FE_OFN328_data_to_iir), 
	.A(data_to_iir));
   CLKBUFX2TS FE_OFC327_data_to_iir (.Y(FE_OFN327_data_to_iir), 
	.A(data_to_iir));
   CLKBUFX2TS FE_OFC326_data_cntl_N191 (.Y(FE_OFN326_data_cntl_N191), 
	.A(\data_cntl/N191 ));
   CLKBUFX2TS FE_OFC325_data_from_fft (.Y(FE_OFN325_data_from_fft), 
	.A(FE_OFN324_data_from_fft));
   CLKBUFX2TS FE_OFC324_data_from_fft (.Y(FE_OFN324_data_from_fft), 
	.A(FE_OFN323_data_from_fft));
   CLKBUFX2TS FE_OFC323_data_from_fft (.Y(FE_OFN323_data_from_fft), 
	.A(data_from_fft));
   CLKBUFX2TS FE_OFC322_data_cntl_N9 (.Y(FE_OFN322_data_cntl_N9), 
	.A(\data_cntl/N9 ));
   CLKBUFX2TS FE_OFC321_data_from_fir (.Y(FE_OFN321_data_from_fir), 
	.A(FE_OFN320_data_from_fir));
   CLKBUFX2TS FE_OFC320_data_from_fir (.Y(FE_OFN320_data_from_fir), 
	.A(FE_OFN319_data_from_fir));
   CLKBUFX2TS FE_OFC319_data_from_fir (.Y(FE_OFN319_data_from_fir), 
	.A(data_from_fir));
   CLKBUFX2TS FE_OFC318_data_cntl_N95 (.Y(FE_OFN318_data_cntl_N95), 
	.A(\data_cntl/N95 ));
   CLKBUFX2TS FE_OFC317_data_from_iir (.Y(FE_OFN317_data_from_iir), 
	.A(FE_OFN316_data_from_iir));
   CLKBUFX2TS FE_OFC316_data_from_iir (.Y(FE_OFN316_data_from_iir), 
	.A(FE_OFN315_data_from_iir));
   CLKBUFX2TS FE_OFC315_data_from_iir (.Y(FE_OFN315_data_from_iir), 
	.A(data_from_iir));
   CLKBUFX2TS FE_OFC314_data_cntl_N159 (.Y(FE_OFN314_data_cntl_N159), 
	.A(\data_cntl/N159 ));
   CLKBUFX2TS FE_OFC313_n2643 (.Y(FE_OFN313_n2643), 
	.A(FE_OFN312_n2643));
   CLKBUFX2TS FE_OFC312_n2643 (.Y(FE_OFN312_n2643), 
	.A(FE_OFN311_n2643));
   CLKBUFX2TS FE_OFC311_n2643 (.Y(FE_OFN311_n2643), 
	.A(FE_OFN310_n2643));
   CLKBUFX3TS FE_OFC310_n2643 (.Y(FE_OFN310_n2643), 
	.A(n2643));
   CLKBUFX2TS FE_OFC309_n2644 (.Y(FE_OFN309_n2644), 
	.A(FE_OFN308_n2644));
   CLKBUFX2TS FE_OFC308_n2644 (.Y(FE_OFN308_n2644), 
	.A(FE_OFN307_n2644));
   CLKBUFX2TS FE_OFC307_n2644 (.Y(FE_OFN307_n2644), 
	.A(FE_OFN306_n2644));
   CLKBUFX3TS FE_OFC306_n2644 (.Y(FE_OFN306_n2644), 
	.A(n2644));
   CLKBUFX2TS FE_OFC305_n2645 (.Y(FE_OFN305_n2645), 
	.A(FE_OFN304_n2645));
   CLKBUFX2TS FE_OFC304_n2645 (.Y(FE_OFN304_n2645), 
	.A(FE_OFN303_n2645));
   CLKBUFX2TS FE_OFC303_n2645 (.Y(FE_OFN303_n2645), 
	.A(FE_OFN302_n2645));
   CLKBUFX3TS FE_OFC302_n2645 (.Y(FE_OFN302_n2645), 
	.A(n2645));
   CLKBUFX2TS FE_OFC301_n2646 (.Y(FE_OFN301_n2646), 
	.A(FE_OFN300_n2646));
   CLKBUFX2TS FE_OFC300_n2646 (.Y(FE_OFN300_n2646), 
	.A(FE_OFN299_n2646));
   CLKBUFX2TS FE_OFC299_n2646 (.Y(FE_OFN299_n2646), 
	.A(FE_OFN298_n2646));
   CLKBUFX3TS FE_OFC298_n2646 (.Y(FE_OFN298_n2646), 
	.A(n2646));
   CLKBUFX2TS FE_OFC297_n2642 (.Y(FE_OFN297_n2642), 
	.A(FE_OFN296_n2642));
   CLKBUFX2TS FE_OFC296_n2642 (.Y(FE_OFN296_n2642), 
	.A(FE_OFN295_n2642));
   CLKBUFX2TS FE_OFC295_n2642 (.Y(FE_OFN295_n2642), 
	.A(FE_OFN294_n2642));
   CLKBUFX3TS FE_OFC294_n2642 (.Y(FE_OFN294_n2642), 
	.A(n2642));
   CLKBUFX2TS FE_OFC293_n2641 (.Y(FE_OFN293_n2641), 
	.A(FE_OFN292_n2641));
   CLKBUFX2TS FE_OFC292_n2641 (.Y(FE_OFN292_n2641), 
	.A(FE_OFN291_n2641));
   CLKBUFX2TS FE_OFC291_n2641 (.Y(FE_OFN291_n2641), 
	.A(FE_OFN289_n2641));
   CLKBUFX2TS FE_OFC290_n2641 (.Y(FE_OFN290_n2641), 
	.A(FE_OFN289_n2641));
   CLKBUFX3TS FE_OFC289_n2641 (.Y(FE_OFN289_n2641), 
	.A(n2641));
   CLKBUFX2TS FE_OFC288_addr_calc_fft_read_calc_count_21_ (.Y(FE_OFN288_addr_calc_fft_read_calc_count_21_), 
	.A(\addr_calc/fft_read_calc/count[21] ));
   BUFX3TS FE_OFC287_addr_calc_fft_read_calc_count_17_ (.Y(FE_OFN287_addr_calc_fft_read_calc_count_17_), 
	.A(\addr_calc/fft_read_calc/count[17] ));
   CLKBUFX2TS FE_OFC286_addr_calc_iir_read_calc_count_30_ (.Y(FE_OFN286_addr_calc_iir_read_calc_count_30_), 
	.A(\addr_calc/iir_read_calc/count[30] ));
   CLKBUFX2TS FE_OFC285_addr_calc_fft_write_calc_count_22_ (.Y(FE_OFN285_addr_calc_fft_write_calc_count_22_), 
	.A(\addr_calc/fft_write_calc/count[22] ));
   CLKBUFX2TS FE_OFC284_addr_calc_fft_write_calc_count_22_ (.Y(FE_OFN284_addr_calc_fft_write_calc_count_22_), 
	.A(\addr_calc/fft_write_calc/count[22] ));
   CLKBUFX2TS FE_OFC283_addr_calc_fir_write_calc_count_20_ (.Y(FE_OFN283_addr_calc_fir_write_calc_count_20_), 
	.A(FE_OFN282_addr_calc_fir_write_calc_count_20_));
   CLKBUFX2TS FE_OFC282_addr_calc_fir_write_calc_count_20_ (.Y(FE_OFN282_addr_calc_fir_write_calc_count_20_), 
	.A(\addr_calc/fir_write_calc/count[20] ));
   CLKBUFX2TS FE_OFC281_addr_calc_fft_write_calc_count_20_ (.Y(FE_OFN281_addr_calc_fft_write_calc_count_20_), 
	.A(FE_OFN280_addr_calc_fft_write_calc_count_20_));
   CLKBUFX2TS FE_OFC280_addr_calc_fft_write_calc_count_20_ (.Y(FE_OFN280_addr_calc_fft_write_calc_count_20_), 
	.A(\addr_calc/fft_write_calc/count[20] ));
   CLKBUFX2TS FE_OFC279_addr_calc_fft_write_calc_count_30_ (.Y(FE_OFN279_addr_calc_fft_write_calc_count_30_), 
	.A(\addr_calc/fft_write_calc/count[30] ));
   CLKBUFX2TS FE_OFC278_addr_calc_fft_read_calc_count_30_ (.Y(FE_OFN278_addr_calc_fft_read_calc_count_30_), 
	.A(\addr_calc/fft_read_calc/count[30] ));
   CLKBUFX2TS FE_OFC277_addr_calc_fft_write_calc_count_24_ (.Y(FE_OFN277_addr_calc_fft_write_calc_count_24_), 
	.A(FE_OFN276_addr_calc_fft_write_calc_count_24_));
   CLKBUFX2TS FE_OFC276_addr_calc_fft_write_calc_count_24_ (.Y(FE_OFN276_addr_calc_fft_write_calc_count_24_), 
	.A(\addr_calc/fft_write_calc/count[24] ));
   CLKBUFX2TS FE_OFC275_addr_calc_fft_read_calc_count_29_ (.Y(FE_OFN275_addr_calc_fft_read_calc_count_29_), 
	.A(\addr_calc/fft_read_calc/count[29] ));
   CLKBUFX2TS FE_OFC274_addr_calc_fft_write_calc_count_31_ (.Y(FE_OFN274_addr_calc_fft_write_calc_count_31_), 
	.A(\addr_calc/fft_write_calc/count[31] ));
   CLKBUFX2TS FE_OFC273_addr_calc_fir_write_calc_count_29_ (.Y(FE_OFN273_addr_calc_fir_write_calc_count_29_), 
	.A(\addr_calc/fir_write_calc/count[29] ));
   CLKBUFX2TS FE_OFC272_addr_calc_fft_write_calc_count_6_ (.Y(FE_OFN272_addr_calc_fft_write_calc_count_6_), 
	.A(\addr_calc/fft_write_calc/count[6] ));
   CLKBUFX2TS FE_OFC271_addr_calc_fft_write_calc_count_6_ (.Y(FE_OFN271_addr_calc_fft_write_calc_count_6_), 
	.A(\addr_calc/fft_write_calc/count[6] ));
   CLKBUFX2TS FE_OFC270_addr_calc_fir_read_calc_count_26_ (.Y(FE_OFN270_addr_calc_fir_read_calc_count_26_), 
	.A(\addr_calc/fir_read_calc/count[26] ));
   CLKBUFX2TS FE_OFC269_addr_calc_fir_read_calc_count_26_ (.Y(FE_OFN269_addr_calc_fir_read_calc_count_26_), 
	.A(\addr_calc/fir_read_calc/count[26] ));
   CLKBUFX2TS FE_OFC268_addr_calc_fir_write_calc_count_26_ (.Y(FE_OFN268_addr_calc_fir_write_calc_count_26_), 
	.A(FE_OFN267_addr_calc_fir_write_calc_count_26_));
   CLKBUFX2TS FE_OFC267_addr_calc_fir_write_calc_count_26_ (.Y(FE_OFN267_addr_calc_fir_write_calc_count_26_), 
	.A(\addr_calc/fir_write_calc/count[26] ));
   CLKBUFX2TS FE_OFC266_addr_calc_iir_write_calc_count_18_ (.Y(FE_OFN266_addr_calc_iir_write_calc_count_18_), 
	.A(\addr_calc/iir_write_calc/count[18] ));
   CLKBUFX2TS FE_OFC265_addr_calc_iir_write_calc_count_18_ (.Y(FE_OFN265_addr_calc_iir_write_calc_count_18_), 
	.A(\addr_calc/iir_write_calc/count[18] ));
   BUFX4TS FE_OFC264_addr_calc_fft_read_calc_count_4_ (.Y(FE_OFN264_addr_calc_fft_read_calc_count_4_), 
	.A(FE_OFN263_addr_calc_fft_read_calc_count_4_));
   CLKBUFX2TS FE_OFC263_addr_calc_fft_read_calc_count_4_ (.Y(FE_OFN263_addr_calc_fft_read_calc_count_4_), 
	.A(\addr_calc/fft_read_calc/count[4] ));
   CLKBUFX2TS FE_OFC262_addr_calc_fir_write_calc_count_31_ (.Y(FE_OFN262_addr_calc_fir_write_calc_count_31_), 
	.A(\addr_calc/fir_write_calc/count[31] ));
   CLKBUFX2TS FE_OFC261_addr_calc_fir_read_calc_count_31_ (.Y(FE_OFN261_addr_calc_fir_read_calc_count_31_), 
	.A(\addr_calc/fir_read_calc/count[31] ));
   BUFX3TS FE_OFC260_addr_calc_fft_write_calc_count_0_ (.Y(FE_OFN260_addr_calc_fft_write_calc_count_0_), 
	.A(\addr_calc/fft_write_calc/count[0] ));
   CLKBUFX2TS FE_OFC259_addr_calc_fft_write_calc_count_14_ (.Y(FE_OFN259_addr_calc_fft_write_calc_count_14_), 
	.A(FE_OFN258_addr_calc_fft_write_calc_count_14_));
   CLKBUFX2TS FE_OFC258_addr_calc_fft_write_calc_count_14_ (.Y(FE_OFN258_addr_calc_fft_write_calc_count_14_), 
	.A(\addr_calc/fft_write_calc/count[14] ));
   BUFX3TS FE_OFC257_addr_calc_fir_write_calc_count_8_ (.Y(FE_OFN257_addr_calc_fir_write_calc_count_8_), 
	.A(FE_OFN256_addr_calc_fir_write_calc_count_8_));
   CLKBUFX2TS FE_OFC256_addr_calc_fir_write_calc_count_8_ (.Y(FE_OFN256_addr_calc_fir_write_calc_count_8_), 
	.A(\addr_calc/fir_write_calc/count[8] ));
   BUFX4TS FE_OFC255_addr_calc_fir_write_calc_count_8_ (.Y(FE_OFN255_addr_calc_fir_write_calc_count_8_), 
	.A(\addr_calc/fir_write_calc/count[8] ));
   CLKBUFX2TS FE_OFC254_addr_calc_fir_write_calc_count_6_ (.Y(FE_OFN254_addr_calc_fir_write_calc_count_6_), 
	.A(FE_OFN253_addr_calc_fir_write_calc_count_6_));
   CLKBUFX2TS FE_OFC253_addr_calc_fir_write_calc_count_6_ (.Y(FE_OFN253_addr_calc_fir_write_calc_count_6_), 
	.A(\addr_calc/fir_write_calc/count[6] ));
   CLKBUFX4TS FE_OFC252_addr_calc_fir_write_calc_count_0_ (.Y(FE_OFN252_addr_calc_fir_write_calc_count_0_), 
	.A(\addr_calc/fir_write_calc/count[0] ));
   CLKBUFX2TS FE_OFC251_addr_calc_fft_read_calc_count_5_ (.Y(FE_OFN251_addr_calc_fft_read_calc_count_5_), 
	.A(\addr_calc/fft_read_calc/count[5] ));
   BUFX6TS FE_OFC250_addr_calc_iir_write_calc_count_3_ (.Y(FE_OFN250_addr_calc_iir_write_calc_count_3_), 
	.A(\addr_calc/iir_write_calc/count[3] ));
   BUFX3TS FE_OFC249_addr_calc_fir_read_calc_count_1_ (.Y(FE_OFN249_addr_calc_fir_read_calc_count_1_), 
	.A(\addr_calc/fir_read_calc/count[1] ));
   CLKBUFX2TS FE_OFC248_addr_calc_iir_read_calc_count_10_ (.Y(FE_OFN248_addr_calc_iir_read_calc_count_10_), 
	.A(\addr_calc/iir_read_calc/count[10] ));
   BUFX3TS FE_OFC247_addr_calc_iir_read_calc_count_7_ (.Y(FE_OFN247_addr_calc_iir_read_calc_count_7_), 
	.A(FE_OFN246_addr_calc_iir_read_calc_count_7_));
   CLKBUFX2TS FE_OFC246_addr_calc_iir_read_calc_count_7_ (.Y(FE_OFN246_addr_calc_iir_read_calc_count_7_), 
	.A(\addr_calc/iir_read_calc/count[7] ));
   CLKBUFX2TS FE_OFC245_addr_calc_fir_read_calc_count_5_ (.Y(FE_OFN245_addr_calc_fir_read_calc_count_5_), 
	.A(\addr_calc/fir_read_calc/count[5] ));
   CLKBUFX2TS FE_OFC244_addr_calc_iir_read_calc_count_4_ (.Y(FE_OFN244_addr_calc_iir_read_calc_count_4_), 
	.A(\addr_calc/iir_read_calc/count[4] ));
   CLKBUFX2TS FE_OFC243_addr_calc_fir_read_calc_count_27_ (.Y(FE_OFN243_addr_calc_fir_read_calc_count_27_), 
	.A(\addr_calc/fir_read_calc/count[27] ));
   CLKBUFX2TS FE_OFC242_addr_calc_fir_write_calc_count_1_ (.Y(FE_OFN242_addr_calc_fir_write_calc_count_1_), 
	.A(\addr_calc/fir_write_calc/count[1] ));
   BUFX12TS FE_OFC241_addr_calc_fir_write_calc_count_4_ (.Y(FE_OFN241_addr_calc_fir_write_calc_count_4_), 
	.A(\addr_calc/fir_write_calc/count[4] ));
   CLKBUFX2TS FE_OFC240_addr_calc_iir_write_calc_count_31_ (.Y(FE_OFN240_addr_calc_iir_write_calc_count_31_), 
	.A(\addr_calc/iir_write_calc/count[31] ));
   CLKBUFX2TS FE_OFC239_addr_calc_iir_write_calc_count_30_ (.Y(FE_OFN239_addr_calc_iir_write_calc_count_30_), 
	.A(\addr_calc/iir_write_calc/count[30] ));
   CLKBUFX2TS FE_OFC238_addr_calc_fir_write_calc_count_30_ (.Y(FE_OFN238_addr_calc_fir_write_calc_count_30_), 
	.A(\addr_calc/fir_write_calc/count[30] ));
   CLKBUFX2TS FE_OFC237_addr_calc_iir_read_calc_count_11_ (.Y(FE_OFN237_addr_calc_iir_read_calc_count_11_), 
	.A(FE_OFN236_addr_calc_iir_read_calc_count_11_));
   CLKBUFX2TS FE_OFC236_addr_calc_iir_read_calc_count_11_ (.Y(FE_OFN236_addr_calc_iir_read_calc_count_11_), 
	.A(\addr_calc/iir_read_calc/count[11] ));
   CLKBUFX2TS FE_OFC235_addr_calc_iir_read_calc_count_27_ (.Y(FE_OFN235_addr_calc_iir_read_calc_count_27_), 
	.A(\addr_calc/iir_read_calc/count[27] ));
   CLKBUFX2TS FE_OFC234_addr_calc_iir_read_calc_count_31_ (.Y(FE_OFN234_addr_calc_iir_read_calc_count_31_), 
	.A(\addr_calc/iir_read_calc/count[31] ));
   CLKBUFX2TS FE_OFC233_addr_calc_fir_write_calc_count_12_ (.Y(FE_OFN233_addr_calc_fir_write_calc_count_12_), 
	.A(\addr_calc/fir_write_calc/count[12] ));
   CLKBUFX2TS FE_OFC232_addr_calc_fir_write_calc_count_12_ (.Y(FE_OFN232_addr_calc_fir_write_calc_count_12_), 
	.A(\addr_calc/fir_write_calc/count[12] ));
   CLKBUFX2TS FE_OFC231_addr_calc_fir_write_calc_count_25_ (.Y(FE_OFN231_addr_calc_fir_write_calc_count_25_), 
	.A(\addr_calc/fir_write_calc/count[25] ));
   CLKBUFX2TS FE_OFC230_addr_calc_iir_write_calc_count_15_ (.Y(FE_OFN230_addr_calc_iir_write_calc_count_15_), 
	.A(FE_OFN229_addr_calc_iir_write_calc_count_15_));
   BUFX3TS FE_OFC229_addr_calc_iir_write_calc_count_15_ (.Y(FE_OFN229_addr_calc_iir_write_calc_count_15_), 
	.A(\addr_calc/iir_write_calc/count[15] ));
   BUFX3TS FE_OFC228_fft_enable (.Y(fft_enable), 
	.A(FE_OFN228_fft_enable));
   CLKBUFX2TS FE_OFC227_addr_calc_fir_read_calc_count_7_ (.Y(FE_OFN227_addr_calc_fir_read_calc_count_7_), 
	.A(\addr_calc/fir_read_calc/count[7] ));
   CLKBUFX2TS FE_OFC226_addr_calc_fft_read_calc_count_31_ (.Y(FE_OFN226_addr_calc_fft_read_calc_count_31_), 
	.A(\addr_calc/fft_read_calc/count[31] ));
   CLKBUFX2TS FE_OFC225_addr_calc_fft_read_calc_count_6_ (.Y(FE_OFN225_addr_calc_fft_read_calc_count_6_), 
	.A(FE_OFN224_addr_calc_fft_read_calc_count_6_));
   CLKBUFX2TS FE_OFC224_addr_calc_fft_read_calc_count_6_ (.Y(FE_OFN224_addr_calc_fft_read_calc_count_6_), 
	.A(\addr_calc/fft_read_calc/count[6] ));
   CLKBUFX2TS FE_OFC223_n643 (.Y(FE_OFN223_n643), 
	.A(FE_OFN222_n643));
   CLKBUFX2TS FE_OFC222_n643 (.Y(FE_OFN222_n643), 
	.A(FE_OFN221_n643));
   CLKBUFX2TS FE_OFC221_n643 (.Y(FE_OFN221_n643), 
	.A(FE_OFN220_n643));
   CLKBUFX2TS FE_OFC220_n643 (.Y(FE_OFN220_n643), 
	.A(FE_OFN219_n643));
   CLKBUFX2TS FE_OFC219_n643 (.Y(FE_OFN219_n643), 
	.A(FE_OFN218_n643));
   CLKBUFX2TS FE_OFC218_n643 (.Y(FE_OFN218_n643), 
	.A(FE_OFN217_n643));
   CLKBUFX2TS FE_OFC217_n643 (.Y(FE_OFN217_n643), 
	.A(FE_OFN216_n643));
   CLKBUFX2TS FE_OFC216_n643 (.Y(FE_OFN216_n643), 
	.A(FE_OFN215_n643));
   CLKBUFX2TS FE_OFC215_n643 (.Y(FE_OFN215_n643), 
	.A(n643));
   CLKBUFX2TS FE_OFC214_n515 (.Y(FE_OFN214_n515), 
	.A(FE_OFN213_n515));
   CLKBUFX2TS FE_OFC213_n515 (.Y(FE_OFN213_n515), 
	.A(FE_OFN211_n515));
   CLKBUFX2TS FE_OFC212_n515 (.Y(FE_OFN212_n515), 
	.A(FE_OFN211_n515));
   CLKBUFX2TS FE_OFC211_n515 (.Y(FE_OFN211_n515), 
	.A(FE_OFN210_n515));
   CLKBUFX2TS FE_OFC210_n515 (.Y(FE_OFN210_n515), 
	.A(FE_OFN209_n515));
   CLKBUFX2TS FE_OFC209_n515 (.Y(FE_OFN209_n515), 
	.A(FE_OFN208_n515));
   CLKBUFX2TS FE_OFC208_n515 (.Y(FE_OFN208_n515), 
	.A(FE_OFN207_n515));
   CLKBUFX2TS FE_OFC207_n515 (.Y(FE_OFN207_n515), 
	.A(n515));
   CLKBUFX2TS FE_OFC206_n387 (.Y(FE_OFN206_n387), 
	.A(FE_OFN204_n387));
   CLKBUFX2TS FE_OFC205_n387 (.Y(FE_OFN205_n387), 
	.A(FE_OFN203_n387));
   CLKBUFX2TS FE_OFC204_n387 (.Y(FE_OFN204_n387), 
	.A(FE_OFN203_n387));
   CLKBUFX2TS FE_OFC203_n387 (.Y(FE_OFN203_n387), 
	.A(FE_OFN202_n387));
   CLKBUFX2TS FE_OFC202_n387 (.Y(FE_OFN202_n387), 
	.A(FE_OFN200_n387));
   CLKBUFX2TS FE_OFC201_n387 (.Y(FE_OFN201_n387), 
	.A(FE_OFN200_n387));
   CLKBUFX2TS FE_OFC200_n387 (.Y(FE_OFN200_n387), 
	.A(FE_OFN198_n387));
   CLKBUFX2TS FE_OFC199_n387 (.Y(FE_OFN199_n387), 
	.A(FE_OFN197_n387));
   CLKBUFX2TS FE_OFC198_n387 (.Y(FE_OFN198_n387), 
	.A(FE_OFN197_n387));
   CLKBUFX2TS FE_OFC197_n387 (.Y(FE_OFN197_n387), 
	.A(n387));
   CLKBUFX2TS FE_OFC196_n707 (.Y(FE_OFN196_n707), 
	.A(FE_OFN195_n707));
   CLKBUFX2TS FE_OFC195_n707 (.Y(FE_OFN195_n707), 
	.A(FE_OFN194_n707));
   CLKBUFX2TS FE_OFC194_n707 (.Y(FE_OFN194_n707), 
	.A(FE_OFN193_n707));
   CLKBUFX2TS FE_OFC193_n707 (.Y(FE_OFN193_n707), 
	.A(FE_OFN192_n707));
   CLKBUFX2TS FE_OFC192_n707 (.Y(FE_OFN192_n707), 
	.A(FE_OFN191_n707));
   CLKBUFX2TS FE_OFC191_n707 (.Y(FE_OFN191_n707), 
	.A(FE_OFN190_n707));
   CLKBUFX2TS FE_OFC190_n707 (.Y(FE_OFN190_n707), 
	.A(n707));
   CLKBUFX2TS FE_OFC189_n579 (.Y(FE_OFN189_n579), 
	.A(FE_OFN188_n579));
   CLKBUFX2TS FE_OFC188_n579 (.Y(FE_OFN188_n579), 
	.A(FE_OFN187_n579));
   CLKBUFX2TS FE_OFC187_n579 (.Y(FE_OFN187_n579), 
	.A(FE_OFN186_n579));
   CLKBUFX2TS FE_OFC186_n579 (.Y(FE_OFN186_n579), 
	.A(FE_OFN185_n579));
   CLKBUFX2TS FE_OFC185_n579 (.Y(FE_OFN185_n579), 
	.A(FE_OFN184_n579));
   CLKBUFX2TS FE_OFC184_n579 (.Y(FE_OFN184_n579), 
	.A(FE_OFN183_n579));
   CLKBUFX2TS FE_OFC183_n579 (.Y(FE_OFN183_n579), 
	.A(n579));
   CLKBUFX2TS FE_OFC182_n451 (.Y(FE_OFN182_n451), 
	.A(FE_OFN181_n451));
   CLKBUFX2TS FE_OFC181_n451 (.Y(FE_OFN181_n451), 
	.A(FE_OFN180_n451));
   CLKBUFX2TS FE_OFC180_n451 (.Y(FE_OFN180_n451), 
	.A(FE_OFN179_n451));
   CLKBUFX2TS FE_OFC179_n451 (.Y(FE_OFN179_n451), 
	.A(FE_OFN178_n451));
   CLKBUFX2TS FE_OFC178_n451 (.Y(FE_OFN178_n451), 
	.A(FE_OFN177_n451));
   CLKBUFX2TS FE_OFC177_n451 (.Y(FE_OFN177_n451), 
	.A(FE_OFN176_n451));
   CLKBUFX2TS FE_OFC176_n451 (.Y(FE_OFN176_n451), 
	.A(n451));
   CLKBUFX2TS FE_OFC175_n131 (.Y(FE_OFN175_n131), 
	.A(FE_OFN174_n131));
   CLKBUFX2TS FE_OFC174_n131 (.Y(FE_OFN174_n131), 
	.A(FE_OFN173_n131));
   CLKBUFX2TS FE_OFC173_n131 (.Y(FE_OFN173_n131), 
	.A(FE_OFN172_n131));
   CLKBUFX2TS FE_OFC172_n131 (.Y(FE_OFN172_n131), 
	.A(n131));
   CLKBUFX2TS FE_OFC171_n195 (.Y(FE_OFN171_n195), 
	.A(FE_OFN170_n195));
   CLKBUFX2TS FE_OFC170_n195 (.Y(FE_OFN170_n195), 
	.A(FE_OFN169_n195));
   CLKBUFX2TS FE_OFC169_n195 (.Y(FE_OFN169_n195), 
	.A(FE_OFN168_n195));
   CLKBUFX2TS FE_OFC168_n195 (.Y(FE_OFN168_n195), 
	.A(n195));
   CLKBUFX2TS FE_OFC167_n259 (.Y(FE_OFN167_n259), 
	.A(FE_OFN166_n259));
   CLKBUFX2TS FE_OFC166_n259 (.Y(FE_OFN166_n259), 
	.A(FE_OFN165_n259));
   CLKBUFX2TS FE_OFC165_n259 (.Y(FE_OFN165_n259), 
	.A(FE_OFN164_n259));
   CLKBUFX2TS FE_OFC164_n259 (.Y(FE_OFN164_n259), 
	.A(n259));
   CLKBUFX2TS FE_OFC163_n323 (.Y(FE_OFN163_n323), 
	.A(FE_OFN162_n323));
   CLKBUFX2TS FE_OFC162_n323 (.Y(FE_OFN162_n323), 
	.A(FE_OFN161_n323));
   CLKBUFX2TS FE_OFC161_n323 (.Y(FE_OFN161_n323), 
	.A(FE_OFN160_n323));
   CLKBUFX2TS FE_OFC160_n323 (.Y(FE_OFN160_n323), 
	.A(n323));
   CLKBUFX2TS FE_OFC159_n67 (.Y(FE_OFN159_n67), 
	.A(FE_OFN158_n67));
   CLKBUFX2TS FE_OFC158_n67 (.Y(FE_OFN158_n67), 
	.A(FE_OFN157_n67));
   CLKBUFX2TS FE_OFC157_n67 (.Y(FE_OFN157_n67), 
	.A(FE_OFN156_n67));
   CLKBUFX2TS FE_OFC156_n67 (.Y(FE_OFN156_n67), 
	.A(n67));
   CLKBUFX2TS FE_OFC155_n3 (.Y(FE_OFN155_n3), 
	.A(FE_OFN154_n3));
   CLKBUFX2TS FE_OFC154_n3 (.Y(FE_OFN154_n3), 
	.A(FE_OFN153_n3));
   CLKBUFX2TS FE_OFC153_n3 (.Y(FE_OFN153_n3), 
	.A(FE_OFN152_n3));
   CLKBUFX2TS FE_OFC152_n3 (.Y(FE_OFN152_n3), 
	.A(n3));
   CLKBUFX2TS FE_OFC151_n2074 (.Y(FE_OFN151_n2074), 
	.A(n2074));
   CLKBUFX2TS FE_OFC150_add_x_22_4_n59 (.Y(FE_OFN150_add_x_22_4_n59), 
	.A(\add_x_22_4/n59 ));
   BUFX3TS FE_OFC149_add_x_22_5_n94 (.Y(FE_OFN149_add_x_22_5_n94), 
	.A(\add_x_22_5/n94 ));
   CLKBUFX2TS FE_OFC148_add_x_22_5_n59 (.Y(FE_OFN148_add_x_22_5_n59), 
	.A(\add_x_22_5/n59 ));
   CLKBUFX2TS FE_OFC147_add_x_22_2_n59 (.Y(FE_OFN147_add_x_22_2_n59), 
	.A(\add_x_22_2/n59 ));
   CLKBUFX2TS FE_OFC146_n801 (.Y(FE_OFN146_n801), 
	.A(FE_OFN145_n801));
   CLKBUFX2TS FE_OFC145_n801 (.Y(FE_OFN145_n801), 
	.A(n801));
   CLKBUFX2TS FE_OFC144_add_x_19_5_n59 (.Y(FE_OFN144_add_x_19_5_n59), 
	.A(\add_x_19_5/n59 ));
   CLKBUFX2TS FE_OFC143_add_x_19_3_n59 (.Y(FE_OFN143_add_x_19_3_n59), 
	.A(\add_x_19_3/n59 ));
   CLKBUFX2TS FE_OFC142_add_x_19_2_n59 (.Y(FE_OFN142_add_x_19_2_n59), 
	.A(\add_x_19_2/n59 ));
   BUFX3TS FE_OFC137_addr_calc_fft_read_addr_10_ (.Y(FE_OFN137_addr_calc_fft_read_addr_10_), 
	.A(\addr_calc/fft_read_addr[10] ));
   CLKBUFX3TS FE_OFC132_addr_calc_fir_write_addr_4_ (.Y(FE_OFN132_addr_calc_fir_write_addr_4_), 
	.A(\addr_calc/fir_write_addr[4] ));
   BUFX6TS FE_OFC131_addr_calc_fir_write_addr_16_ (.Y(FE_OFN131_addr_calc_fir_write_addr_16_), 
	.A(\addr_calc/fir_write_addr[16] ));
   BUFX16TS FE_OFC129_add_x_19_5_n157 (.Y(FE_OFN129_add_x_19_5_n157), 
	.A(\add_x_19_5/n157 ));
   BUFX12TS FE_OFC122_add_x_19_2_n157 (.Y(FE_OFN122_add_x_19_2_n157), 
	.A(\add_x_19_2/n157 ));
   BUFX3TS FE_OFC121_addr_calc_iir_read_addr_4_ (.Y(FE_OFN121_addr_calc_iir_read_addr_4_), 
	.A(\addr_calc/iir_read_addr[4] ));
   BUFX6TS FE_OFC117_addr_calc_iir_read_addr_10_ (.Y(FE_OFN117_addr_calc_iir_read_addr_10_), 
	.A(\addr_calc/iir_read_addr[10] ));
   BUFX3TS FE_OFC114_DP_OP_159_297_3515_n852 (.Y(FE_OFN114_DP_OP_159_297_3515_n852), 
	.A(\DP_OP_159_297_3515/n852 ));
   CLKBUFX2TS FE_OFC93_n1192 (.Y(FE_OFN93_n1192), 
	.A(FE_OFN92_n1192));
   CLKBUFX2TS FE_OFC92_n1192 (.Y(FE_OFN92_n1192), 
	.A(FE_OFN91_n1192));
   CLKBUFX2TS FE_OFC91_n1192 (.Y(FE_OFN91_n1192), 
	.A(FE_OFN90_n1192));
   BUFX3TS FE_OFC90_n1192 (.Y(FE_OFN90_n1192), 
	.A(n1192));
   CLKBUFX2TS FE_OFC89_n2654 (.Y(FE_OFN89_n2654), 
	.A(FE_OFN88_n2654));
   CLKBUFX2TS FE_OFC88_n2654 (.Y(FE_OFN88_n2654), 
	.A(FE_OFN87_n2654));
   CLKBUFX2TS FE_OFC87_n2654 (.Y(FE_OFN87_n2654), 
	.A(FE_OFN86_n2654));
   BUFX3TS FE_OFC86_n2654 (.Y(FE_OFN86_n2654), 
	.A(FE_OFN85_n2654));
   BUFX3TS FE_OFC85_n2654 (.Y(FE_OFN85_n2654), 
	.A(n2654));
   CLKBUFX3TS FE_OFC84_n2787 (.Y(FE_OFN84_n2787), 
	.A(FE_OFN83_n2787));
   BUFX3TS FE_OFC83_n2787 (.Y(FE_OFN83_n2787), 
	.A(FE_OFN82_n2787));
   BUFX3TS FE_OFC82_n2787 (.Y(FE_OFN82_n2787), 
	.A(FE_OFN81_n2787));
   BUFX3TS FE_OFC81_n2787 (.Y(FE_OFN81_n2787), 
	.A(FE_OFN80_n2787));
   BUFX3TS FE_OFC80_n2787 (.Y(FE_OFN80_n2787), 
	.A(FE_OFN79_n2787));
   BUFX8TS FE_OFC79_n2787 (.Y(FE_OFN79_n2787), 
	.A(FE_OFN78_n2787));
   BUFX3TS FE_OFC78_n2787 (.Y(FE_OFN78_n2787), 
	.A(FE_OCPUNCON1880_n2787));
   BUFX6TS FE_OFC75_n2599 (.Y(FE_OFN75_n2599), 
	.A(n2599));
   BUFX3TS FE_OFC71_n2809 (.Y(FE_OFN71_n2809), 
	.A(FE_OFN70_n2809));
   BUFX3TS FE_OFC70_n2809 (.Y(FE_OFN70_n2809), 
	.A(FE_OFN69_n2809));
   BUFX3TS FE_OFC69_n2809 (.Y(FE_OFN69_n2809), 
	.A(FE_OFN68_n2809));
   BUFX3TS FE_OFC68_n2809 (.Y(FE_OFN68_n2809), 
	.A(FE_OFN67_n2809));
   BUFX3TS FE_OFC67_n2809 (.Y(FE_OFN67_n2809), 
	.A(FE_OFN66_n2809));
   BUFX3TS FE_OFC66_n2809 (.Y(FE_OFN66_n2809), 
	.A(FE_OFN65_n2809));
   BUFX3TS FE_OFC65_n2809 (.Y(FE_OFN65_n2809), 
	.A(FE_OFN64_n2809));
   BUFX3TS FE_OFC64_n2809 (.Y(FE_OFN64_n2809), 
	.A(FE_OFN63_n2809));
   BUFX3TS FE_OFC63_n2809 (.Y(FE_OFN63_n2809), 
	.A(FE_OFN62_n2809));
   BUFX3TS FE_OFC62_n2809 (.Y(FE_OFN62_n2809), 
	.A(n2809));
   BUFX3TS FE_OFC61_n2807 (.Y(FE_OFN61_n2807), 
	.A(FE_OFN60_n2807));
   BUFX3TS FE_OFC60_n2807 (.Y(FE_OFN60_n2807), 
	.A(FE_OFN59_n2807));
   BUFX3TS FE_OFC59_n2807 (.Y(FE_OFN59_n2807), 
	.A(FE_OFN58_n2807));
   BUFX3TS FE_OFC58_n2807 (.Y(FE_OFN58_n2807), 
	.A(FE_OFN57_n2807));
   BUFX3TS FE_OFC57_n2807 (.Y(FE_OFN57_n2807), 
	.A(FE_OFN56_n2807));
   BUFX3TS FE_OFC56_n2807 (.Y(FE_OFN56_n2807), 
	.A(FE_OFN55_n2807));
   BUFX3TS FE_OFC55_n2807 (.Y(FE_OFN55_n2807), 
	.A(FE_OFN53_n2807));
   CLKBUFX2TS FE_OFC54_n2807 (.Y(FE_OFN54_n2807), 
	.A(FE_OFN53_n2807));
   BUFX3TS FE_OFC53_n2807 (.Y(FE_OFN53_n2807), 
	.A(FE_OFN52_n2807));
   BUFX3TS FE_OFC52_n2807 (.Y(FE_OFN52_n2807), 
	.A(n2807));
   BUFX4TS FE_OFC51_n2803 (.Y(FE_OFN51_n2803), 
	.A(FE_OFN50_n2803));
   BUFX4TS FE_OFC50_n2803 (.Y(FE_OFN50_n2803), 
	.A(FE_OFN49_n2803));
   BUFX8TS FE_OFC49_n2803 (.Y(FE_OFN49_n2803), 
	.A(FE_OFN48_n2803));
   BUFX3TS FE_OFC48_n2803 (.Y(FE_OFN48_n2803), 
	.A(FE_OFN547_n2803));
   BUFX16TS FE_OFC47_n1758 (.Y(FE_OFN47_n1758), 
	.A(n1758));
   BUFX20TS FE_OFC35_n2795 (.Y(FE_OFN35_n2795), 
	.A(FE_OFN34_n2795));
   BUFX8TS FE_OFC34_n2795 (.Y(FE_OFN34_n2795), 
	.A(FE_OFN33_n2795));
   BUFX3TS FE_OFC33_n2795 (.Y(FE_OFN33_n2795), 
	.A(FE_OFN32_n2795));
   BUFX3TS FE_OFC32_n2795 (.Y(FE_OFN32_n2795), 
	.A(FE_OFN31_n2795));
   BUFX20TS FE_OFC31_n2795 (.Y(FE_OFN31_n2795), 
	.A(FE_OFN30_n2795));
   BUFX8TS FE_OFC30_n2795 (.Y(FE_OFN30_n2795), 
	.A(FE_OFN29_n2795));
   BUFX3TS FE_OFC29_n2795 (.Y(FE_OFN29_n2795), 
	.A(FE_OFN28_n2795));
   BUFX8TS FE_OFC28_n2795 (.Y(FE_OFN28_n2795), 
	.A(FE_OFN27_n2795));
   BUFX3TS FE_OFC27_n2795 (.Y(FE_OFN27_n2795), 
	.A(n2795));
   BUFX3TS FE_OFC26_n2797 (.Y(FE_OFN26_n2797), 
	.A(FE_OFN25_n2797));
   BUFX8TS FE_OFC25_n2797 (.Y(FE_OFN25_n2797), 
	.A(FE_OFN24_n2797));
   BUFX3TS FE_OFC24_n2797 (.Y(FE_OFN24_n2797), 
	.A(FE_OFN23_n2797));
   BUFX3TS FE_OFC23_n2797 (.Y(FE_OFN23_n2797), 
	.A(FE_OFN22_n2797));
   BUFX3TS FE_OFC22_n2797 (.Y(FE_OFN22_n2797), 
	.A(FE_OFN21_n2797));
   BUFX3TS FE_OFC21_n2797 (.Y(FE_OFN21_n2797), 
	.A(FE_OFN20_n2797));
   BUFX3TS FE_OFC20_n2797 (.Y(FE_OFN20_n2797), 
	.A(FE_OFN19_n2797));
   BUFX8TS FE_OFC19_n2797 (.Y(FE_OFN19_n2797), 
	.A(FE_OFN18_n2797));
   BUFX3TS FE_OFC18_n2797 (.Y(FE_OFN18_n2797), 
	.A(FE_OFN17_n2797));
   BUFX8TS FE_OFC17_n2797 (.Y(FE_OFN17_n2797), 
	.A(n2797));
   BUFX3TS FE_OFC16_n2794 (.Y(FE_OFN16_n2794), 
	.A(FE_OFN15_n2794));
   BUFX3TS FE_OFC15_n2794 (.Y(FE_OFN15_n2794), 
	.A(FE_OFN14_n2794));
   BUFX3TS FE_OFC14_n2794 (.Y(FE_OFN14_n2794), 
	.A(FE_OFN13_n2794));
   BUFX3TS FE_OFC13_n2794 (.Y(FE_OFN13_n2794), 
	.A(FE_OFN12_n2794));
   BUFX3TS FE_OFC12_n2794 (.Y(FE_OFN12_n2794), 
	.A(FE_OFN11_n2794));
   BUFX3TS FE_OFC11_n2794 (.Y(FE_OFN11_n2794), 
	.A(FE_OFN10_n2794));
   BUFX3TS FE_OFC10_n2794 (.Y(FE_OFN10_n2794), 
	.A(FE_OFN9_n2794));
   BUFX3TS FE_OFC9_n2794 (.Y(FE_OFN9_n2794), 
	.A(FE_OFN8_n2794));
   BUFX3TS FE_OFC8_n2794 (.Y(FE_OFN8_n2794), 
	.A(FE_OFN7_n2794));
   BUFX3TS FE_OFC7_n2794 (.Y(FE_OFN7_n2794), 
	.A(n2794));
   CLKBUFX2TS FE_OFC6_n1750 (.Y(FE_OFN6_n1750), 
	.A(FE_OFN552_n1751));
   CLKBUFX2TS FE_OFC4_n1755 (.Y(FE_OFN4_n1755), 
	.A(n1755));
   BUFX3TS FE_OFC3_n1754 (.Y(FE_OFN3_n1754), 
	.A(FE_OFN2_n1754));
   CLKBUFX3TS FE_OFC2_n1754 (.Y(FE_OFN2_n1754), 
	.A(n1754));
   CLKBUFX2TS FE_OFC1_n1751 (.Y(FE_OFN1_n1751), 
	.A(FE_OFN552_n1751));
   NOR4X1TS U71 (.Y(n816), 
	.D(n2580), 
	.C(FE_OFN248_addr_calc_iir_read_calc_count_10_), 
	.B(FE_OFN236_addr_calc_iir_read_calc_count_11_), 
	.A(n1785));
   NOR4X1TS U197 (.Y(n846), 
	.D(n1924), 
	.C(n2020), 
	.B(\addr_calc/fft_write_calc/count[19] ), 
	.A(n1941));
   NOR4X1TS U274 (.Y(n867), 
	.D(\addr_calc/fir_write_calc/count[0] ), 
	.C(\addr_calc/fir_write_calc/count[10] ), 
	.B(n1877), 
	.A(FE_OFN233_addr_calc_fir_write_calc_count_12_));
   NOR4X1TS U288 (.Y(n883), 
	.D(\addr_calc/fir_read_calc/count[13] ), 
	.C(\addr_calc/fir_read_calc/count[14] ), 
	.B(\addr_calc/fir_read_calc/count[15] ), 
	.A(\addr_calc/fir_read_calc/count[16] ));
   NOR4X1TS U289 (.Y(n882), 
	.D(n2007), 
	.C(\addr_calc/fir_read_calc/count[10] ), 
	.B(n1895), 
	.A(n1994));
   NOR4X1TS U291 (.Y(n880), 
	.D(\addr_calc/fir_read_calc/count[17] ), 
	.C(n1988), 
	.B(\addr_calc/fir_read_calc/count[19] ), 
	.A(\addr_calc/fir_read_calc/count[1] ));
   NAND3X1TS U294 (.Y(n885), 
	.C(n886), 
	.B(n2066), 
	.A(FE_OFN145_n801));
   NAND3BX1TS U299 (.Y(n897), 
	.C(fir_read_done), 
	.B(fir_write_done), 
	.AN(n884));
   OAI33XLTS U306 (.Y(n1135), 
	.B2(iir_write_done), 
	.B1(n869), 
	.B0(n899), 
	.A2(n1861), 
	.A1(n901), 
	.A0(n891));
   NAND2X1TS U310 (.Y(n870), 
	.B(n2311), 
	.A(n902));
   NAND2X1TS U313 (.Y(n899), 
	.B(n872), 
	.A(FE_OFN335_instruction_2_));
   NAND3X1TS U315 (.Y(n903), 
	.C(n906), 
	.B(n905), 
	.A(n904));
   NAND3BX1TS U323 (.Y(n907), 
	.C(\pla_top/instruction_valid ), 
	.B(FE_OFN336_instruction_0_), 
	.AN(instruction[9]));
   NOR4X1TS U338 (.Y(n921), 
	.D(n2578), 
	.C(n1940), 
	.B(n1942), 
	.A(n2044));
   OA21X2TS U343 (.Y(iir_get_req), 
	.B0(iir_get_req_reg), 
	.A1(n923), 
	.A0(n796));
   OA21X2TS U350 (.Y(fir_get_req), 
	.B0(fir_get_req_reg), 
	.A1(n927), 
	.A0(n798));
   NOR4XLTS U365 (.Y(\data_cntl/N256 ), 
	.D(n932), 
	.C(n933), 
	.B(FE_OFN516_from_iir_full), 
	.A(FE_OFN514_to_iir_full));
   NOR4XLTS U371 (.Y(\data_cntl/N253 ), 
	.D(n1830), 
	.C(n937), 
	.B(FE_OFN512_from_fir_full), 
	.A(FE_OFN510_to_fir_full));
   NAND3X1TS U381 (.Y(n932), 
	.C(FE_OFN560_n2587), 
	.B(FE_OFN563_n2060), 
	.A(n2815));
   TLATXLTS \data_cntl/fft_get_req_reg  (.QN(n929), 
	.G(\data_cntl/N260 ), 
	.D(\data_cntl/N261 ));
   TLATXLTS \data_cntl/fft_put_req_reg  (.Q(fft_put_req_reg), 
	.G(\data_cntl/N260 ), 
	.D(\data_cntl/N259 ));
   TLATXLTS \data_cntl/fir_put_req_reg  (.Q(fir_put_req_reg), 
	.G(\data_cntl/N263 ), 
	.D(\data_cntl/N262 ));
   TLATXLTS \data_cntl/iir_put_req_reg  (.Q(iir_put_req_reg), 
	.G(\data_cntl/N266 ), 
	.D(\data_cntl/N265 ));
   TLATXLTS \data_cntl/iir_get_req_reg  (.Q(iir_get_req_reg), 
	.G(\data_cntl/N266 ), 
	.D(\data_cntl/N267 ));
   TLATXLTS \data_cntl/fir_get_req_reg  (.Q(fir_get_req_reg), 
	.G(\data_cntl/N263 ), 
	.D(\data_cntl/N264 ));
   TLATXLTS \data_cntl/data_to_fft_reg  (.QN(\data_cntl/N63 ), 
	.Q(data_to_fft), 
	.G(\data_cntl/N250 ), 
	.D(\data_cntl/N251 ));
   TLATXLTS \data_cntl/data_to_fir_reg  (.QN(\data_cntl/N99 ), 
	.Q(data_to_fir), 
	.G(\data_cntl/N255 ), 
	.D(\data_cntl/N253 ));
   TLATXLTS \data_cntl/data_to_iir_reg  (.QN(\data_cntl/N191 ), 
	.Q(data_to_iir), 
	.G(\data_cntl/N258 ), 
	.D(\data_cntl/N256 ));
   TLATXLTS \data_cntl/data_from_fft_reg  (.QN(\data_cntl/N9 ), 
	.Q(data_from_fft), 
	.G(\data_cntl/N250 ), 
	.D(\data_cntl/N252 ));
   TLATXLTS \data_cntl/data_from_fir_reg  (.QN(\data_cntl/N95 ), 
	.Q(data_from_fir), 
	.G(\data_cntl/N255 ), 
	.D(\data_cntl/N254 ));
   TLATXLTS \data_cntl/data_from_iir_reg  (.QN(\data_cntl/N159 ), 
	.Q(data_from_iir), 
	.G(\data_cntl/N258 ), 
	.D(\data_cntl/N257 ));
   TLATXLTS \addr_calc/from_fir_go_reg  (.QN(\addr_calc/N99 ), 
	.Q(n2643), 
	.G(\addr_calc/N220 ), 
	.D(\data_cntl/N264 ));
   TLATXLTS \addr_calc/to_fir_go_reg  (.QN(\addr_calc/N95 ), 
	.Q(n2644), 
	.G(\addr_calc/N220 ), 
	.D(\addr_calc/N219 ));
   TLATXLTS \addr_calc/from_fft_go_reg  (.QN(\addr_calc/N63 ), 
	.Q(n2645), 
	.G(\addr_calc/N216 ), 
	.D(\data_cntl/N261 ));
   TLATXLTS \addr_calc/to_fft_go_reg  (.QN(\addr_calc/N9 ), 
	.Q(n2646), 
	.G(\addr_calc/N216 ), 
	.D(\addr_calc/N217 ));
   TLATXLTS \addr_calc/to_iir_go_reg  (.QN(\addr_calc/N159 ), 
	.Q(n2642), 
	.G(\addr_calc/N224 ), 
	.D(\addr_calc/N223 ));
   TLATXLTS \addr_calc/from_iir_go_reg  (.QN(\addr_calc/N191 ), 
	.Q(n2641), 
	.G(\addr_calc/N224 ), 
	.D(\data_cntl/N267 ));
   DFFQX4TS \pla_top/acc_done_reg  (.Q(acc_done), 
	.D(n1134), 
	.CK(clk__L1_N0));
   TBUFX2TS \data_cntl/fft_data_out_tri[31]  (.Y(fft_data_out[31]), 
	.OE(FE_OFN334_data_to_fft), 
	.A(n2360));
   TBUFX2TS \data_cntl/fft_data_out_tri[30]  (.Y(fft_data_out[30]), 
	.OE(FE_OFN334_data_to_fft), 
	.A(n2502));
   TBUFX2TS \data_cntl/fft_data_out_tri[29]  (.Y(fft_data_out[29]), 
	.OE(FE_OFN334_data_to_fft), 
	.A(n2518));
   TBUFX2TS \data_cntl/fft_data_out_tri[28]  (.Y(fft_data_out[28]), 
	.OE(FE_OFN334_data_to_fft), 
	.A(n2534));
   TBUFX2TS \data_cntl/fft_data_out_tri[27]  (.Y(fft_data_out[27]), 
	.OE(FE_OFN215_n643), 
	.A(n2356));
   TBUFX2TS \data_cntl/fft_data_out_tri[26]  (.Y(fft_data_out[26]), 
	.OE(n643), 
	.A(n2504));
   TBUFX2TS \data_cntl/fft_data_out_tri[25]  (.Y(fft_data_out[25]), 
	.OE(FE_OFN215_n643), 
	.A(n2520));
   TBUFX2TS \data_cntl/fft_data_out_tri[24]  (.Y(fft_data_out[24]), 
	.OE(FE_OFN215_n643), 
	.A(n2536));
   TBUFX2TS \data_cntl/fft_data_out_tri[23]  (.Y(fft_data_out[23]), 
	.OE(FE_OFN216_n643), 
	.A(n2352));
   TBUFX2TS \data_cntl/fft_data_out_tri[22]  (.Y(fft_data_out[22]), 
	.OE(FE_OFN217_n643), 
	.A(n2506));
   TBUFX2TS \data_cntl/fft_data_out_tri[21]  (.Y(fft_data_out[21]), 
	.OE(FE_OFN220_n643), 
	.A(n2522));
   TBUFX2TS \data_cntl/fft_data_out_tri[20]  (.Y(fft_data_out[20]), 
	.OE(FE_OFN221_n643), 
	.A(n2538));
   TBUFX2TS \data_cntl/fft_data_out_tri[19]  (.Y(fft_data_out[19]), 
	.OE(FE_OFN218_n643), 
	.A(n2348));
   TBUFX2TS \data_cntl/fft_data_out_tri[18]  (.Y(fft_data_out[18]), 
	.OE(FE_OFN219_n643), 
	.A(n2508));
   TBUFX2TS \data_cntl/fft_data_out_tri[17]  (.Y(fft_data_out[17]), 
	.OE(FE_OFN217_n643), 
	.A(n2524));
   TBUFX2TS \data_cntl/fft_data_out_tri[16]  (.Y(fft_data_out[16]), 
	.OE(FE_OFN222_n643), 
	.A(n2540));
   TBUFX2TS \data_cntl/fft_data_out_tri[15]  (.Y(fft_data_out[15]), 
	.OE(FE_OFN219_n643), 
	.A(n2346));
   TBUFX2TS \data_cntl/fft_data_out_tri[14]  (.Y(fft_data_out[14]), 
	.OE(FE_OFN223_n643), 
	.A(n2510));
   TBUFX2TS \data_cntl/fft_data_out_tri[13]  (.Y(fft_data_out[13]), 
	.OE(FE_OFN221_n643), 
	.A(n2526));
   TBUFX2TS \data_cntl/fft_data_out_tri[12]  (.Y(fft_data_out[12]), 
	.OE(FE_OFN216_n643), 
	.A(n2542));
   TBUFX2TS \data_cntl/fft_data_out_tri[11]  (.Y(fft_data_out[11]), 
	.OE(FE_OFN217_n643), 
	.A(n2350));
   TBUFX2TS \data_cntl/fft_data_out_tri[10]  (.Y(fft_data_out[10]), 
	.OE(FE_OFN216_n643), 
	.A(n2512));
   TBUFX2TS \data_cntl/fft_data_out_tri[9]  (.Y(fft_data_out[9]), 
	.OE(FE_OFN222_n643), 
	.A(n2528));
   TBUFX2TS \data_cntl/fft_data_out_tri[8]  (.Y(fft_data_out[8]), 
	.OE(FE_OFN222_n643), 
	.A(n2544));
   TBUFX2TS \data_cntl/fft_data_out_tri[7]  (.Y(fft_data_out[7]), 
	.OE(FE_OFN221_n643), 
	.A(n2354));
   TBUFX2TS \data_cntl/fft_data_out_tri[6]  (.Y(fft_data_out[6]), 
	.OE(FE_OFN219_n643), 
	.A(n2514));
   TBUFX2TS \data_cntl/fft_data_out_tri[5]  (.Y(fft_data_out[5]), 
	.OE(FE_OFN220_n643), 
	.A(n2530));
   TBUFX2TS \data_cntl/fft_data_out_tri[4]  (.Y(fft_data_out[4]), 
	.OE(FE_OFN223_n643), 
	.A(n2546));
   TBUFX2TS \data_cntl/fft_data_out_tri[3]  (.Y(fft_data_out[3]), 
	.OE(FE_OFN218_n643), 
	.A(n2358));
   TBUFX2TS \data_cntl/fft_data_out_tri[2]  (.Y(fft_data_out[2]), 
	.OE(FE_OFN223_n643), 
	.A(n2516));
   TBUFX2TS \data_cntl/fft_data_out_tri[1]  (.Y(fft_data_out[1]), 
	.OE(FE_OFN223_n643), 
	.A(n2532));
   TBUFX2TS \data_cntl/fft_data_out_tri[0]  (.Y(fft_data_out[0]), 
	.OE(FE_OFN220_n643), 
	.A(n2548));
   TBUFX2TS \data_cntl/fir_data_out_tri[31]  (.Y(fir_data_out[31]), 
	.OE(FE_OFN331_data_to_fir), 
	.A(n2360));
   TBUFX2TS \data_cntl/fir_data_out_tri[30]  (.Y(fir_data_out[30]), 
	.OE(FE_OFN331_data_to_fir), 
	.A(n2502));
   TBUFX2TS \data_cntl/fir_data_out_tri[29]  (.Y(fir_data_out[29]), 
	.OE(FE_OFN331_data_to_fir), 
	.A(n2518));
   TBUFX2TS \data_cntl/fir_data_out_tri[28]  (.Y(fir_data_out[28]), 
	.OE(FE_OFN331_data_to_fir), 
	.A(n2534));
   TBUFX2TS \data_cntl/fir_data_out_tri[27]  (.Y(fir_data_out[27]), 
	.OE(n515), 
	.A(n2356));
   TBUFX2TS \data_cntl/fir_data_out_tri[26]  (.Y(fir_data_out[26]), 
	.OE(n515), 
	.A(n2504));
   TBUFX2TS \data_cntl/fir_data_out_tri[25]  (.Y(fir_data_out[25]), 
	.OE(n515), 
	.A(n2520));
   TBUFX2TS \data_cntl/fir_data_out_tri[24]  (.Y(fir_data_out[24]), 
	.OE(FE_OFN207_n515), 
	.A(n2536));
   TBUFX2TS \data_cntl/fir_data_out_tri[23]  (.Y(fir_data_out[23]), 
	.OE(FE_OFN210_n515), 
	.A(n2352));
   TBUFX2TS \data_cntl/fir_data_out_tri[22]  (.Y(fir_data_out[22]), 
	.OE(FE_OFN208_n515), 
	.A(n2506));
   TBUFX2TS \data_cntl/fir_data_out_tri[21]  (.Y(fir_data_out[21]), 
	.OE(FE_OFN211_n515), 
	.A(n2522));
   TBUFX2TS \data_cntl/fir_data_out_tri[20]  (.Y(fir_data_out[20]), 
	.OE(FE_OFN214_n515), 
	.A(n2538));
   TBUFX2TS \data_cntl/fir_data_out_tri[19]  (.Y(fir_data_out[19]), 
	.OE(FE_OFN209_n515), 
	.A(n2348));
   TBUFX2TS \data_cntl/fir_data_out_tri[18]  (.Y(fir_data_out[18]), 
	.OE(FE_OFN212_n515), 
	.A(n2508));
   TBUFX2TS \data_cntl/fir_data_out_tri[17]  (.Y(fir_data_out[17]), 
	.OE(FE_OFN208_n515), 
	.A(n2524));
   TBUFX2TS \data_cntl/fir_data_out_tri[16]  (.Y(fir_data_out[16]), 
	.OE(FE_OFN211_n515), 
	.A(n2540));
   TBUFX2TS \data_cntl/fir_data_out_tri[15]  (.Y(fir_data_out[15]), 
	.OE(FE_OFN212_n515), 
	.A(n2346));
   TBUFX2TS \data_cntl/fir_data_out_tri[14]  (.Y(fir_data_out[14]), 
	.OE(FE_OFN213_n515), 
	.A(n2510));
   TBUFX2TS \data_cntl/fir_data_out_tri[13]  (.Y(fir_data_out[13]), 
	.OE(FE_OFN212_n515), 
	.A(n2526));
   TBUFX2TS \data_cntl/fir_data_out_tri[12]  (.Y(fir_data_out[12]), 
	.OE(FE_OFN207_n515), 
	.A(n2542));
   TBUFX2TS \data_cntl/fir_data_out_tri[11]  (.Y(fir_data_out[11]), 
	.OE(FE_OFN209_n515), 
	.A(n2350));
   TBUFX2TS \data_cntl/fir_data_out_tri[10]  (.Y(fir_data_out[10]), 
	.OE(FE_OFN207_n515), 
	.A(n2512));
   TBUFX2TS \data_cntl/fir_data_out_tri[9]  (.Y(fir_data_out[9]), 
	.OE(FE_OFN210_n515), 
	.A(n2528));
   TBUFX2TS \data_cntl/fir_data_out_tri[8]  (.Y(fir_data_out[8]), 
	.OE(FE_OFN214_n515), 
	.A(n2544));
   TBUFX2TS \data_cntl/fir_data_out_tri[7]  (.Y(fir_data_out[7]), 
	.OE(FE_OFN212_n515), 
	.A(n2354));
   TBUFX2TS \data_cntl/fir_data_out_tri[6]  (.Y(fir_data_out[6]), 
	.OE(FE_OFN209_n515), 
	.A(n2514));
   TBUFX2TS \data_cntl/fir_data_out_tri[5]  (.Y(fir_data_out[5]), 
	.OE(FE_OFN213_n515), 
	.A(n2530));
   TBUFX2TS \data_cntl/fir_data_out_tri[4]  (.Y(fir_data_out[4]), 
	.OE(FE_OFN213_n515), 
	.A(n2546));
   TBUFX2TS \data_cntl/fir_data_out_tri[3]  (.Y(fir_data_out[3]), 
	.OE(FE_OFN208_n515), 
	.A(n2358));
   TBUFX2TS \data_cntl/fir_data_out_tri[2]  (.Y(fir_data_out[2]), 
	.OE(FE_OFN214_n515), 
	.A(n2516));
   TBUFX2TS \data_cntl/fir_data_out_tri[1]  (.Y(fir_data_out[1]), 
	.OE(FE_OFN214_n515), 
	.A(n2532));
   TBUFX2TS \data_cntl/fir_data_out_tri[0]  (.Y(fir_data_out[0]), 
	.OE(FE_OFN210_n515), 
	.A(n2548));
   TBUFX2TS \data_cntl/iir_data_out_tri[31]  (.Y(iir_data_out[31]), 
	.OE(FE_OFN328_data_to_iir), 
	.A(n2360));
   TBUFX2TS \data_cntl/iir_data_out_tri[30]  (.Y(iir_data_out[30]), 
	.OE(FE_OFN328_data_to_iir), 
	.A(n2502));
   TBUFX2TS \data_cntl/iir_data_out_tri[29]  (.Y(iir_data_out[29]), 
	.OE(FE_OFN328_data_to_iir), 
	.A(n2518));
   TBUFX2TS \data_cntl/iir_data_out_tri[28]  (.Y(iir_data_out[28]), 
	.OE(FE_OFN328_data_to_iir), 
	.A(n2534));
   TBUFX2TS \data_cntl/iir_data_out_tri[27]  (.Y(iir_data_out[27]), 
	.OE(FE_OFN199_n387), 
	.A(n2356));
   TBUFX2TS \data_cntl/iir_data_out_tri[26]  (.Y(iir_data_out[26]), 
	.OE(FE_OFN199_n387), 
	.A(n2504));
   TBUFX2TS \data_cntl/iir_data_out_tri[25]  (.Y(iir_data_out[25]), 
	.OE(FE_OFN197_n387), 
	.A(n2520));
   TBUFX2TS \data_cntl/iir_data_out_tri[24]  (.Y(iir_data_out[24]), 
	.OE(FE_OFN199_n387), 
	.A(n2536));
   TBUFX2TS \data_cntl/iir_data_out_tri[23]  (.Y(iir_data_out[23]), 
	.OE(FE_OFN201_n387), 
	.A(n2352));
   TBUFX2TS \data_cntl/iir_data_out_tri[22]  (.Y(iir_data_out[22]), 
	.OE(FE_OFN198_n387), 
	.A(n2506));
   TBUFX2TS \data_cntl/iir_data_out_tri[21]  (.Y(iir_data_out[21]), 
	.OE(FE_OFN203_n387), 
	.A(n2522));
   TBUFX2TS \data_cntl/iir_data_out_tri[20]  (.Y(iir_data_out[20]), 
	.OE(FE_OFN205_n387), 
	.A(n2538));
   TBUFX2TS \data_cntl/iir_data_out_tri[19]  (.Y(iir_data_out[19]), 
	.OE(FE_OFN198_n387), 
	.A(n2348));
   TBUFX2TS \data_cntl/iir_data_out_tri[18]  (.Y(iir_data_out[18]), 
	.OE(FE_OFN205_n387), 
	.A(n2508));
   TBUFX2TS \data_cntl/iir_data_out_tri[17]  (.Y(iir_data_out[17]), 
	.OE(n387), 
	.A(n2524));
   TBUFX2TS \data_cntl/iir_data_out_tri[16]  (.Y(iir_data_out[16]), 
	.OE(FE_OFN204_n387), 
	.A(n2540));
   TBUFX2TS \data_cntl/iir_data_out_tri[15]  (.Y(iir_data_out[15]), 
	.OE(FE_OFN202_n387), 
	.A(n2346));
   TBUFX2TS \data_cntl/iir_data_out_tri[14]  (.Y(iir_data_out[14]), 
	.OE(FE_OFN206_n387), 
	.A(n2510));
   TBUFX2TS \data_cntl/iir_data_out_tri[13]  (.Y(iir_data_out[13]), 
	.OE(FE_OFN205_n387), 
	.A(n2526));
   TBUFX2TS \data_cntl/iir_data_out_tri[12]  (.Y(iir_data_out[12]), 
	.OE(FE_OFN199_n387), 
	.A(n2542));
   TBUFX2TS \data_cntl/iir_data_out_tri[11]  (.Y(iir_data_out[11]), 
	.OE(FE_OFN201_n387), 
	.A(n2350));
   TBUFX2TS \data_cntl/iir_data_out_tri[10]  (.Y(iir_data_out[10]), 
	.OE(FE_OFN197_n387), 
	.A(n2512));
   TBUFX2TS \data_cntl/iir_data_out_tri[9]  (.Y(iir_data_out[9]), 
	.OE(FE_OFN204_n387), 
	.A(n2528));
   TBUFX2TS \data_cntl/iir_data_out_tri[8]  (.Y(iir_data_out[8]), 
	.OE(FE_OFN203_n387), 
	.A(n2544));
   TBUFX2TS \data_cntl/iir_data_out_tri[7]  (.Y(iir_data_out[7]), 
	.OE(FE_OFN205_n387), 
	.A(n2354));
   TBUFX2TS \data_cntl/iir_data_out_tri[6]  (.Y(iir_data_out[6]), 
	.OE(FE_OFN200_n387), 
	.A(n2514));
   TBUFX2TS \data_cntl/iir_data_out_tri[5]  (.Y(iir_data_out[5]), 
	.OE(FE_OFN202_n387), 
	.A(n2530));
   TBUFX2TS \data_cntl/iir_data_out_tri[4]  (.Y(iir_data_out[4]), 
	.OE(n387), 
	.A(n2546));
   TBUFX2TS \data_cntl/iir_data_out_tri[3]  (.Y(iir_data_out[3]), 
	.OE(FE_OFN200_n387), 
	.A(n2358));
   TBUFX2TS \data_cntl/iir_data_out_tri[2]  (.Y(iir_data_out[2]), 
	.OE(FE_OFN206_n387), 
	.A(n2516));
   TBUFX2TS \data_cntl/iir_data_out_tri[1]  (.Y(iir_data_out[1]), 
	.OE(FE_OFN206_n387), 
	.A(n2532));
   TBUFX2TS \data_cntl/iir_data_out_tri[0]  (.Y(iir_data_out[0]), 
	.OE(FE_OFN202_n387), 
	.A(n2548));
   TBUFX2TS \data_cntl/data_bus_tri[31]  (.Y(data_bus[31]), 
	.OE(FE_OFN324_data_from_fft), 
	.A(fft_data_in[31]));
   TBUFX2TS \data_cntl/data_bus_tri[30]  (.Y(data_bus[30]), 
	.OE(FE_OFN323_data_from_fft), 
	.A(fft_data_in[30]));
   TBUFX2TS \data_cntl/data_bus_tri[29]  (.Y(data_bus[29]), 
	.OE(FE_OFN324_data_from_fft), 
	.A(fft_data_in[29]));
   TBUFX2TS \data_cntl/data_bus_tri[28]  (.Y(data_bus[28]), 
	.OE(FE_OFN324_data_from_fft), 
	.A(fft_data_in[28]));
   TBUFX2TS \data_cntl/data_bus_tri[27]  (.Y(data_bus[27]), 
	.OE(FE_OFN325_data_from_fft), 
	.A(fft_data_in[27]));
   TBUFX2TS \data_cntl/data_bus_tri[26]  (.Y(data_bus[26]), 
	.OE(FE_OFN325_data_from_fft), 
	.A(fft_data_in[26]));
   TBUFX2TS \data_cntl/data_bus_tri[25]  (.Y(data_bus[25]), 
	.OE(FE_OFN325_data_from_fft), 
	.A(fft_data_in[25]));
   TBUFX2TS \data_cntl/data_bus_tri[24]  (.Y(data_bus[24]), 
	.OE(FE_OFN325_data_from_fft), 
	.A(fft_data_in[24]));
   TBUFX2TS \data_cntl/data_bus_tri[23]  (.Y(data_bus[23]), 
	.OE(FE_OFN191_n707), 
	.A(fft_data_in[23]));
   TBUFX2TS \data_cntl/data_bus_tri[22]  (.Y(data_bus[22]), 
	.OE(FE_OFN194_n707), 
	.A(fft_data_in[22]));
   TBUFX2TS \data_cntl/data_bus_tri[21]  (.Y(data_bus[21]), 
	.OE(FE_OFN196_n707), 
	.A(fft_data_in[21]));
   TBUFX2TS \data_cntl/data_bus_tri[20]  (.Y(data_bus[20]), 
	.OE(FE_OFN194_n707), 
	.A(fft_data_in[20]));
   TBUFX2TS \data_cntl/data_bus_tri[19]  (.Y(data_bus[19]), 
	.OE(FE_OFN196_n707), 
	.A(fft_data_in[19]));
   TBUFX2TS \data_cntl/data_bus_tri[18]  (.Y(data_bus[18]), 
	.OE(FE_OFN190_n707), 
	.A(fft_data_in[18]));
   TBUFX2TS \data_cntl/data_bus_tri[17]  (.Y(data_bus[17]), 
	.OE(FE_OFN192_n707), 
	.A(fft_data_in[17]));
   TBUFX2TS \data_cntl/data_bus_tri[16]  (.Y(data_bus[16]), 
	.OE(FE_OFN192_n707), 
	.A(fft_data_in[16]));
   TBUFX2TS \data_cntl/data_bus_tri[15]  (.Y(data_bus[15]), 
	.OE(FE_OFN192_n707), 
	.A(fft_data_in[15]));
   TBUFX2TS \data_cntl/data_bus_tri[14]  (.Y(data_bus[14]), 
	.OE(FE_OFN191_n707), 
	.A(fft_data_in[14]));
   TBUFX2TS \data_cntl/data_bus_tri[13]  (.Y(data_bus[13]), 
	.OE(FE_OFN196_n707), 
	.A(fft_data_in[13]));
   TBUFX2TS \data_cntl/data_bus_tri[12]  (.Y(data_bus[12]), 
	.OE(n707), 
	.A(fft_data_in[12]));
   TBUFX2TS \data_cntl/data_bus_tri[11]  (.Y(data_bus[11]), 
	.OE(FE_OFN193_n707), 
	.A(fft_data_in[11]));
   TBUFX2TS \data_cntl/data_bus_tri[10]  (.Y(data_bus[10]), 
	.OE(n707), 
	.A(fft_data_in[10]));
   TBUFX2TS \data_cntl/data_bus_tri[9]  (.Y(data_bus[9]), 
	.OE(FE_OFN194_n707), 
	.A(FE_OFN503_fft_data_in_9_));
   TBUFX2TS \data_cntl/data_bus_tri[8]  (.Y(data_bus[8]), 
	.OE(FE_OFN191_n707), 
	.A(fft_data_in[8]));
   TBUFX2TS \data_cntl/data_bus_tri[7]  (.Y(data_bus[7]), 
	.OE(FE_OFN190_n707), 
	.A(fft_data_in[7]));
   TBUFX2TS \data_cntl/data_bus_tri[6]  (.Y(data_bus[6]), 
	.OE(FE_OFN193_n707), 
	.A(fft_data_in[6]));
   TBUFX2TS \data_cntl/data_bus_tri[5]  (.Y(data_bus[5]), 
	.OE(FE_OFN196_n707), 
	.A(fft_data_in[5]));
   TBUFX2TS \data_cntl/data_bus_tri[4]  (.Y(data_bus[4]), 
	.OE(FE_OFN195_n707), 
	.A(fft_data_in[4]));
   TBUFX2TS \data_cntl/data_bus_tri[3]  (.Y(data_bus[3]), 
	.OE(FE_OFN195_n707), 
	.A(fft_data_in[3]));
   TBUFX2TS \data_cntl/data_bus_tri[2]  (.Y(data_bus[2]), 
	.OE(FE_OFN193_n707), 
	.A(fft_data_in[2]));
   TBUFX2TS \data_cntl/data_bus_tri[1]  (.Y(data_bus[1]), 
	.OE(FE_OFN195_n707), 
	.A(fft_data_in[1]));
   TBUFX2TS \data_cntl/data_bus_tri[0]  (.Y(data_bus[0]), 
	.OE(FE_OFN190_n707), 
	.A(fft_data_in[0]));
   TBUFX2TS \data_cntl/data_bus_tri2[31]  (.Y(data_bus[31]), 
	.OE(FE_OFN320_data_from_fir), 
	.A(fir_data_in[31]));
   TBUFX2TS \data_cntl/data_bus_tri2[30]  (.Y(data_bus[30]), 
	.OE(FE_OFN319_data_from_fir), 
	.A(fir_data_in[30]));
   TBUFX2TS \data_cntl/data_bus_tri2[29]  (.Y(data_bus[29]), 
	.OE(FE_OFN321_data_from_fir), 
	.A(fir_data_in[29]));
   TBUFX2TS \data_cntl/data_bus_tri2[28]  (.Y(data_bus[28]), 
	.OE(FE_OFN320_data_from_fir), 
	.A(fir_data_in[28]));
   TBUFX2TS \data_cntl/data_bus_tri2[27]  (.Y(data_bus[27]), 
	.OE(FE_OFN320_data_from_fir), 
	.A(fir_data_in[27]));
   TBUFX2TS \data_cntl/data_bus_tri2[26]  (.Y(data_bus[26]), 
	.OE(FE_OFN321_data_from_fir), 
	.A(fir_data_in[26]));
   TBUFX2TS \data_cntl/data_bus_tri2[25]  (.Y(data_bus[25]), 
	.OE(FE_OFN321_data_from_fir), 
	.A(fir_data_in[25]));
   TBUFX2TS \data_cntl/data_bus_tri2[24]  (.Y(data_bus[24]), 
	.OE(FE_OFN321_data_from_fir), 
	.A(fir_data_in[24]));
   TBUFX2TS \data_cntl/data_bus_tri2[23]  (.Y(data_bus[23]), 
	.OE(FE_OFN184_n579), 
	.A(fir_data_in[23]));
   TBUFX2TS \data_cntl/data_bus_tri2[22]  (.Y(data_bus[22]), 
	.OE(FE_OFN188_n579), 
	.A(fir_data_in[22]));
   TBUFX2TS \data_cntl/data_bus_tri2[21]  (.Y(data_bus[21]), 
	.OE(FE_OFN189_n579), 
	.A(fir_data_in[21]));
   TBUFX2TS \data_cntl/data_bus_tri2[20]  (.Y(data_bus[20]), 
	.OE(FE_OFN187_n579), 
	.A(fir_data_in[20]));
   TBUFX2TS \data_cntl/data_bus_tri2[19]  (.Y(data_bus[19]), 
	.OE(FE_OFN189_n579), 
	.A(fir_data_in[19]));
   TBUFX2TS \data_cntl/data_bus_tri2[18]  (.Y(data_bus[18]), 
	.OE(FE_OFN183_n579), 
	.A(fir_data_in[18]));
   TBUFX2TS \data_cntl/data_bus_tri2[17]  (.Y(data_bus[17]), 
	.OE(FE_OFN184_n579), 
	.A(fir_data_in[17]));
   TBUFX2TS \data_cntl/data_bus_tri2[16]  (.Y(data_bus[16]), 
	.OE(FE_OFN185_n579), 
	.A(fir_data_in[16]));
   TBUFX2TS \data_cntl/data_bus_tri2[15]  (.Y(data_bus[15]), 
	.OE(FE_OFN185_n579), 
	.A(fir_data_in[15]));
   TBUFX2TS \data_cntl/data_bus_tri2[14]  (.Y(data_bus[14]), 
	.OE(FE_OFN185_n579), 
	.A(fir_data_in[14]));
   TBUFX2TS \data_cntl/data_bus_tri2[13]  (.Y(data_bus[13]), 
	.OE(FE_OFN188_n579), 
	.A(fir_data_in[13]));
   TBUFX2TS \data_cntl/data_bus_tri2[12]  (.Y(data_bus[12]), 
	.OE(n579), 
	.A(fir_data_in[12]));
   TBUFX2TS \data_cntl/data_bus_tri2[11]  (.Y(data_bus[11]), 
	.OE(FE_OFN186_n579), 
	.A(fir_data_in[11]));
   TBUFX2TS \data_cntl/data_bus_tri2[10]  (.Y(data_bus[10]), 
	.OE(n579), 
	.A(fir_data_in[10]));
   TBUFX2TS \data_cntl/data_bus_tri2[9]  (.Y(data_bus[9]), 
	.OE(FE_OFN187_n579), 
	.A(fir_data_in[9]));
   TBUFX2TS \data_cntl/data_bus_tri2[8]  (.Y(data_bus[8]), 
	.OE(FE_OFN183_n579), 
	.A(fir_data_in[8]));
   TBUFX2TS \data_cntl/data_bus_tri2[7]  (.Y(data_bus[7]), 
	.OE(FE_OFN184_n579), 
	.A(fir_data_in[7]));
   TBUFX2TS \data_cntl/data_bus_tri2[6]  (.Y(data_bus[6]), 
	.OE(FE_OFN187_n579), 
	.A(fir_data_in[6]));
   TBUFX2TS \data_cntl/data_bus_tri2[5]  (.Y(data_bus[5]), 
	.OE(FE_OFN189_n579), 
	.A(fir_data_in[5]));
   TBUFX2TS \data_cntl/data_bus_tri2[4]  (.Y(data_bus[4]), 
	.OE(FE_OFN188_n579), 
	.A(fir_data_in[4]));
   TBUFX2TS \data_cntl/data_bus_tri2[3]  (.Y(data_bus[3]), 
	.OE(FE_OFN186_n579), 
	.A(fir_data_in[3]));
   TBUFX2TS \data_cntl/data_bus_tri2[2]  (.Y(data_bus[2]), 
	.OE(FE_OFN186_n579), 
	.A(fir_data_in[2]));
   TBUFX2TS \data_cntl/data_bus_tri2[1]  (.Y(data_bus[1]), 
	.OE(FE_OFN189_n579), 
	.A(fir_data_in[1]));
   TBUFX2TS \data_cntl/data_bus_tri2[0]  (.Y(data_bus[0]), 
	.OE(FE_OFN183_n579), 
	.A(fir_data_in[0]));
   TBUFX2TS \data_cntl/data_bus_tri3[31]  (.Y(data_bus[31]), 
	.OE(FE_OFN317_data_from_iir), 
	.A(iir_data_in[31]));
   TBUFX2TS \data_cntl/data_bus_tri3[30]  (.Y(data_bus[30]), 
	.OE(FE_OFN317_data_from_iir), 
	.A(iir_data_in[30]));
   TBUFX2TS \data_cntl/data_bus_tri3[29]  (.Y(data_bus[29]), 
	.OE(FE_OFN317_data_from_iir), 
	.A(iir_data_in[29]));
   TBUFX2TS \data_cntl/data_bus_tri3[28]  (.Y(data_bus[28]), 
	.OE(FE_OFN317_data_from_iir), 
	.A(iir_data_in[28]));
   TBUFX2TS \data_cntl/data_bus_tri3[27]  (.Y(data_bus[27]), 
	.OE(FE_OFN316_data_from_iir), 
	.A(iir_data_in[27]));
   TBUFX2TS \data_cntl/data_bus_tri3[26]  (.Y(data_bus[26]), 
	.OE(FE_OFN315_data_from_iir), 
	.A(iir_data_in[26]));
   TBUFX2TS \data_cntl/data_bus_tri3[25]  (.Y(data_bus[25]), 
	.OE(FE_OFN316_data_from_iir), 
	.A(iir_data_in[25]));
   TBUFX2TS \data_cntl/data_bus_tri3[24]  (.Y(data_bus[24]), 
	.OE(FE_OFN316_data_from_iir), 
	.A(iir_data_in[24]));
   TBUFX2TS \data_cntl/data_bus_tri3[23]  (.Y(data_bus[23]), 
	.OE(FE_OFN177_n451), 
	.A(iir_data_in[23]));
   TBUFX2TS \data_cntl/data_bus_tri3[22]  (.Y(data_bus[22]), 
	.OE(FE_OFN181_n451), 
	.A(iir_data_in[22]));
   TBUFX2TS \data_cntl/data_bus_tri3[21]  (.Y(data_bus[21]), 
	.OE(FE_OFN182_n451), 
	.A(iir_data_in[21]));
   TBUFX2TS \data_cntl/data_bus_tri3[20]  (.Y(data_bus[20]), 
	.OE(FE_OFN179_n451), 
	.A(iir_data_in[20]));
   TBUFX2TS \data_cntl/data_bus_tri3[19]  (.Y(data_bus[19]), 
	.OE(FE_OFN182_n451), 
	.A(iir_data_in[19]));
   TBUFX2TS \data_cntl/data_bus_tri3[18]  (.Y(data_bus[18]), 
	.OE(FE_OFN176_n451), 
	.A(iir_data_in[18]));
   TBUFX2TS \data_cntl/data_bus_tri3[17]  (.Y(data_bus[17]), 
	.OE(FE_OFN178_n451), 
	.A(iir_data_in[17]));
   TBUFX2TS \data_cntl/data_bus_tri3[16]  (.Y(data_bus[16]), 
	.OE(FE_OFN178_n451), 
	.A(iir_data_in[16]));
   TBUFX2TS \data_cntl/data_bus_tri3[15]  (.Y(data_bus[15]), 
	.OE(FE_OFN178_n451), 
	.A(iir_data_in[15]));
   TBUFX2TS \data_cntl/data_bus_tri3[14]  (.Y(data_bus[14]), 
	.OE(FE_OFN177_n451), 
	.A(iir_data_in[14]));
   TBUFX2TS \data_cntl/data_bus_tri3[13]  (.Y(data_bus[13]), 
	.OE(FE_OFN182_n451), 
	.A(iir_data_in[13]));
   TBUFX2TS \data_cntl/data_bus_tri3[12]  (.Y(data_bus[12]), 
	.OE(n451), 
	.A(iir_data_in[12]));
   TBUFX2TS \data_cntl/data_bus_tri3[11]  (.Y(data_bus[11]), 
	.OE(FE_OFN179_n451), 
	.A(iir_data_in[11]));
   TBUFX2TS \data_cntl/data_bus_tri3[10]  (.Y(data_bus[10]), 
	.OE(n451), 
	.A(iir_data_in[10]));
   TBUFX2TS \data_cntl/data_bus_tri3[9]  (.Y(data_bus[9]), 
	.OE(FE_OFN180_n451), 
	.A(FE_OFN504_iir_data_in_9_));
   TBUFX2TS \data_cntl/data_bus_tri3[8]  (.Y(data_bus[8]), 
	.OE(FE_OFN176_n451), 
	.A(iir_data_in[8]));
   TBUFX2TS \data_cntl/data_bus_tri3[7]  (.Y(data_bus[7]), 
	.OE(FE_OFN177_n451), 
	.A(iir_data_in[7]));
   TBUFX2TS \data_cntl/data_bus_tri3[6]  (.Y(data_bus[6]), 
	.OE(FE_OFN180_n451), 
	.A(iir_data_in[6]));
   TBUFX2TS \data_cntl/data_bus_tri3[5]  (.Y(data_bus[5]), 
	.OE(FE_OFN182_n451), 
	.A(iir_data_in[5]));
   TBUFX2TS \data_cntl/data_bus_tri3[4]  (.Y(data_bus[4]), 
	.OE(FE_OFN181_n451), 
	.A(iir_data_in[4]));
   TBUFX2TS \data_cntl/data_bus_tri3[3]  (.Y(data_bus[3]), 
	.OE(FE_OFN180_n451), 
	.A(iir_data_in[3]));
   TBUFX2TS \data_cntl/data_bus_tri3[2]  (.Y(data_bus[2]), 
	.OE(FE_OFN179_n451), 
	.A(iir_data_in[2]));
   TBUFX2TS \data_cntl/data_bus_tri3[1]  (.Y(data_bus[1]), 
	.OE(FE_OFN181_n451), 
	.A(iir_data_in[1]));
   TBUFX2TS \data_cntl/data_bus_tri3[0]  (.Y(data_bus[0]), 
	.OE(FE_OFN176_n451), 
	.A(iir_data_in[0]));
   TBUFX3TS \addr_calc/addr_tri[0]  (.Y(addr[0]), 
	.OE(FE_OFN301_n2646), 
	.A(\addr_calc/fft_read_addr[0] ));
   TBUFX3TS \addr_calc/addr_tri2[0]  (.Y(addr[0]), 
	.OE(FE_OFN305_n2645), 
	.A(\addr_calc/fft_write_addr[0] ));
   TBUFX3TS \addr_calc/addr_tri3[0]  (.Y(addr[0]), 
	.OE(FE_OFN309_n2644), 
	.A(\addr_calc/fir_read_addr[0] ));
   TBUFX3TS \addr_calc/addr_tri4[0]  (.Y(addr[0]), 
	.OE(FE_OFN313_n2643), 
	.A(\addr_calc/fir_write_addr[0] ));
   TBUFX3TS \addr_calc/addr_tri5[0]  (.Y(addr[0]), 
	.OE(FE_OFN297_n2642), 
	.A(\addr_calc/iir_read_addr[0] ));
   TBUFX3TS \addr_calc/addr_tri6[0]  (.Y(addr[0]), 
	.OE(FE_OFN293_n2641), 
	.A(\addr_calc/iir_write_addr[0] ));
   TBUFX2TS \addr_calc/addr_tri[3]  (.Y(addr[3]), 
	.OE(FE_OFN301_n2646), 
	.A(\addr_calc/fft_read_addr[3] ));
   TBUFX2TS \addr_calc/addr_tri2[4]  (.Y(addr[4]), 
	.OE(FE_OFN167_n259), 
	.A(\addr_calc/fft_write_addr[4] ));
   TBUFX2TS \addr_calc/addr_tri2[3]  (.Y(addr[3]), 
	.OE(FE_OFN305_n2645), 
	.A(\addr_calc/fft_write_addr[3] ));
   TBUFX2TS \addr_calc/addr_tri3[4]  (.Y(addr[4]), 
	.OE(FE_OFN171_n195), 
	.A(\addr_calc/fir_read_addr[4] ));
   TBUFX2TS \addr_calc/addr_tri3[3]  (.Y(addr[3]), 
	.OE(FE_OFN309_n2644), 
	.A(\addr_calc/fir_read_addr[3] ));
   TBUFX2TS \addr_calc/addr_tri4[4]  (.Y(addr[4]), 
	.OE(FE_OFN175_n131), 
	.A(FE_OFN132_addr_calc_fir_write_addr_4_));
   TBUFX2TS \addr_calc/addr_tri4[3]  (.Y(addr[3]), 
	.OE(FE_OFN313_n2643), 
	.A(\addr_calc/fir_write_addr[3] ));
   TBUFX2TS \addr_calc/addr_tri5[3]  (.Y(addr[3]), 
	.OE(FE_OFN297_n2642), 
	.A(\addr_calc/iir_read_addr[3] ));
   TBUFX2TS \addr_calc/addr_tri6[4]  (.Y(addr[4]), 
	.OE(FE_OFN155_n3), 
	.A(\addr_calc/iir_write_addr[4] ));
   TBUFX3TS \addr_calc/addr_tri6[3]  (.Y(addr[3]), 
	.OE(FE_OFN293_n2641), 
	.A(\addr_calc/iir_write_addr[3] ));
   TBUFX3TS \addr_calc/addr_tri[1]  (.Y(addr[1]), 
	.OE(FE_OFN301_n2646), 
	.A(\addr_calc/fft_read_addr[1] ));
   TBUFX2TS \addr_calc/addr_tri2[2]  (.Y(addr[2]), 
	.OE(FE_OFN305_n2645), 
	.A(\addr_calc/fft_write_addr[2] ));
   TBUFX3TS \addr_calc/addr_tri2[1]  (.Y(addr[1]), 
	.OE(FE_OFN305_n2645), 
	.A(\addr_calc/fft_write_addr[1] ));
   TBUFX2TS \addr_calc/addr_tri3[2]  (.Y(addr[2]), 
	.OE(FE_OFN309_n2644), 
	.A(\addr_calc/fir_read_addr[2] ));
   TBUFX3TS \addr_calc/addr_tri3[1]  (.Y(addr[1]), 
	.OE(FE_OFN309_n2644), 
	.A(\addr_calc/fir_read_addr[1] ));
   TBUFX2TS \addr_calc/addr_tri4[2]  (.Y(addr[2]), 
	.OE(FE_OFN313_n2643), 
	.A(\addr_calc/fir_write_addr[2] ));
   TBUFX3TS \addr_calc/addr_tri4[1]  (.Y(addr[1]), 
	.OE(FE_OFN313_n2643), 
	.A(\addr_calc/fir_write_addr[1] ));
   TBUFX3TS \addr_calc/addr_tri5[1]  (.Y(addr[1]), 
	.OE(FE_OFN297_n2642), 
	.A(\addr_calc/iir_read_addr[1] ));
   TBUFX2TS \addr_calc/addr_tri6[2]  (.Y(addr[2]), 
	.OE(FE_OFN293_n2641), 
	.A(\addr_calc/iir_write_addr[2] ));
   TBUFX3TS \addr_calc/addr_tri6[1]  (.Y(addr[1]), 
	.OE(FE_OFN293_n2641), 
	.A(\addr_calc/iir_write_addr[1] ));
   DFFQX1TS \pla_top/instruction_valid_reg  (.Q(\pla_top/instruction_valid ), 
	.D(\pla_top/N59 ), 
	.CK(clk__L1_N0));
   DFFQX4TS \pla_top/iir_enable_reg  (.Q(n2815), 
	.D(n1135), 
	.CK(clk__L1_N0));
   TBUFX16TS \addr_calc/addr_tri[29]  (.Y(addr[29]), 
	.OE(FE_OFN300_n2646), 
	.A(FE_OFN136_addr_calc_fft_read_addr_29_));
   TBUFX3TS \addr_calc/addr_tri[16]  (.Y(addr[16]), 
	.OE(FE_OFN160_n323), 
	.A(\addr_calc/fft_read_addr[16] ));
   TBUFX4TS \addr_calc/addr_tri[13]  (.Y(addr[13]), 
	.OE(n323), 
	.A(\addr_calc/fft_read_addr[13] ));
   TBUFX3TS \addr_calc/addr_tri[10]  (.Y(addr[10]), 
	.OE(n2646), 
	.A(FE_OFN137_addr_calc_fft_read_addr_10_));
   TBUFX4TS \addr_calc/addr_tri[9]  (.Y(addr[9]), 
	.OE(n2646), 
	.A(\addr_calc/fft_read_addr[9] ));
   TBUFX2TS \addr_calc/addr_tri[7]  (.Y(addr[7]), 
	.OE(FE_OFN163_n323), 
	.A(FE_OFN532_addr_calc_fft_read_addr_7_));
   TBUFX2TS \addr_calc/addr_tri[4]  (.Y(addr[4]), 
	.OE(FE_OFN163_n323), 
	.A(\addr_calc/fft_read_addr[4] ));
   TBUFX16TS \addr_calc/addr_tri2[29]  (.Y(addr[29]), 
	.OE(FE_OFN304_n2645), 
	.A(\addr_calc/fft_write_addr[29] ));
   TBUFX2TS \addr_calc/addr_tri2[16]  (.Y(addr[16]), 
	.OE(FE_OFN164_n259), 
	.A(\addr_calc/fft_write_addr[16] ));
   TBUFX2TS \addr_calc/addr_tri2[10]  (.Y(addr[10]), 
	.OE(n2645), 
	.A(\addr_calc/fft_write_addr[10] ));
   TBUFX3TS \addr_calc/addr_tri2[9]  (.Y(addr[9]), 
	.OE(n2645), 
	.A(\addr_calc/fft_write_addr[9] ));
   TBUFX2TS \addr_calc/addr_tri2[7]  (.Y(addr[7]), 
	.OE(FE_OFN167_n259), 
	.A(\addr_calc/fft_write_addr[7] ));
   TBUFX8TS \addr_calc/addr_tri3[29]  (.Y(addr[29]), 
	.OE(FE_OFN308_n2644), 
	.A(\addr_calc/fir_read_addr[29] ));
   TBUFX2TS \addr_calc/addr_tri3[16]  (.Y(addr[16]), 
	.OE(FE_OFN168_n195), 
	.A(\addr_calc/fir_read_addr[16] ));
   TBUFX3TS \addr_calc/addr_tri3[10]  (.Y(addr[10]), 
	.OE(n2644), 
	.A(\addr_calc/fir_read_addr[10] ));
   TBUFX4TS \addr_calc/addr_tri3[9]  (.Y(addr[9]), 
	.OE(n2644), 
	.A(\addr_calc/fir_read_addr[9] ));
   TBUFX2TS \addr_calc/addr_tri3[7]  (.Y(addr[7]), 
	.OE(FE_OFN171_n195), 
	.A(\addr_calc/fir_read_addr[7] ));
   TBUFX16TS \addr_calc/addr_tri4[29]  (.Y(addr[29]), 
	.OE(FE_OFN312_n2643), 
	.A(\addr_calc/fir_write_addr[29] ));
   TBUFX8TS \addr_calc/addr_tri4[16]  (.Y(addr[16]), 
	.OE(FE_OFN172_n131), 
	.A(FE_OFN131_addr_calc_fir_write_addr_16_));
   TBUFX2TS \addr_calc/addr_tri4[10]  (.Y(addr[10]), 
	.OE(n2643), 
	.A(\addr_calc/fir_write_addr[10] ));
   TBUFX2TS \addr_calc/addr_tri4[9]  (.Y(addr[9]), 
	.OE(n2643), 
	.A(\addr_calc/fir_write_addr[9] ));
   TBUFX2TS \addr_calc/addr_tri4[7]  (.Y(addr[7]), 
	.OE(FE_OFN175_n131), 
	.A(FE_OFN533_addr_calc_fir_write_addr_7_));
   TBUFX6TS \addr_calc/addr_tri5[16]  (.Y(addr[16]), 
	.OE(FE_OFN156_n67), 
	.A(\addr_calc/iir_read_addr[16] ));
   TBUFX3TS \addr_calc/addr_tri5[10]  (.Y(addr[10]), 
	.OE(n2642), 
	.A(FE_OFN117_addr_calc_iir_read_addr_10_));
   TBUFX3TS \addr_calc/addr_tri5[9]  (.Y(addr[9]), 
	.OE(n2642), 
	.A(FE_OFN541_addr_calc_iir_read_addr_9_));
   TBUFX8TS \addr_calc/addr_tri5[7]  (.Y(addr[7]), 
	.OE(FE_OFN159_n67), 
	.A(FE_OFN536_addr_calc_iir_read_addr_7_));
   TBUFX2TS \addr_calc/addr_tri5[4]  (.Y(addr[4]), 
	.OE(FE_OFN159_n67), 
	.A(FE_OFN121_addr_calc_iir_read_addr_4_));
   TBUFX12TS \addr_calc/addr_tri6[29]  (.Y(addr[29]), 
	.OE(FE_OFN292_n2641), 
	.A(\addr_calc/iir_write_addr[29] ));
   TBUFX2TS \addr_calc/addr_tri6[16]  (.Y(addr[16]), 
	.OE(FE_OFN152_n3), 
	.A(FE_OFN124_addr_calc_iir_write_addr_16_));
   TBUFX2TS \addr_calc/addr_tri6[10]  (.Y(addr[10]), 
	.OE(FE_OFN290_n2641), 
	.A(FE_OFN128_addr_calc_iir_write_addr_10_));
   TBUFX2TS \addr_calc/addr_tri6[9]  (.Y(addr[9]), 
	.OE(FE_OFN290_n2641), 
	.A(FE_OFN127_addr_calc_iir_write_addr_9_));
   TBUFX2TS \addr_calc/addr_tri6[7]  (.Y(addr[7]), 
	.OE(FE_OFN155_n3), 
	.A(FE_OFN534_addr_calc_iir_write_addr_7_));
   TBUFX16TS \addr_calc/addr_tri[12]  (.Y(addr[12]), 
	.OE(n323), 
	.A(\addr_calc/fft_read_addr[12] ));
   TBUFX4TS \addr_calc/addr_tri[11]  (.Y(addr[11]), 
	.OE(n2646), 
	.A(FE_OFN544_addr_calc_fft_read_addr_11_));
   TBUFX4TS \addr_calc/addr_tri[8]  (.Y(addr[8]), 
	.OE(FE_OFN298_n2646), 
	.A(\addr_calc/fft_read_addr[8] ));
   TBUFX2TS \addr_calc/addr_tri[6]  (.Y(addr[6]), 
	.OE(FE_OFN163_n323), 
	.A(\addr_calc/fft_read_addr[6] ));
   TBUFX2TS \addr_calc/addr_tri[5]  (.Y(addr[5]), 
	.OE(FE_OFN163_n323), 
	.A(\addr_calc/fft_read_addr[5] ));
   TBUFX2TS \addr_calc/addr_tri[2]  (.Y(addr[2]), 
	.OE(FE_OFN301_n2646), 
	.A(\addr_calc/fft_read_addr[2] ));
   TBUFX3TS \addr_calc/addr_tri2[24]  (.Y(addr[24]), 
	.OE(FE_OFN302_n2645), 
	.A(\addr_calc/fft_write_addr[24] ));
   TBUFX16TS \addr_calc/addr_tri2[20]  (.Y(addr[20]), 
	.OE(FE_OFN165_n259), 
	.A(\addr_calc/fft_write_addr[20] ));
   TBUFX8TS \addr_calc/addr_tri2[12]  (.Y(addr[12]), 
	.OE(n259), 
	.A(\addr_calc/fft_write_addr[12] ));
   TBUFX2TS \addr_calc/addr_tri2[11]  (.Y(addr[11]), 
	.OE(n2645), 
	.A(\addr_calc/fft_write_addr[11] ));
   TBUFX2TS \addr_calc/addr_tri2[8]  (.Y(addr[8]), 
	.OE(FE_OFN302_n2645), 
	.A(\addr_calc/fft_write_addr[8] ));
   TBUFX2TS \addr_calc/addr_tri2[6]  (.Y(addr[6]), 
	.OE(FE_OFN167_n259), 
	.A(\addr_calc/fft_write_addr[6] ));
   TBUFX2TS \addr_calc/addr_tri2[5]  (.Y(addr[5]), 
	.OE(FE_OFN167_n259), 
	.A(\addr_calc/fft_write_addr[5] ));
   TBUFX8TS \addr_calc/addr_tri3[24]  (.Y(addr[24]), 
	.OE(FE_OFN306_n2644), 
	.A(\addr_calc/fir_read_addr[24] ));
   TBUFX4TS \addr_calc/addr_tri3[14]  (.Y(addr[14]), 
	.OE(n195), 
	.A(\addr_calc/fir_read_addr[14] ));
   TBUFX2TS \addr_calc/addr_tri3[12]  (.Y(addr[12]), 
	.OE(n195), 
	.A(\addr_calc/fir_read_addr[12] ));
   TBUFX8TS \addr_calc/addr_tri3[11]  (.Y(addr[11]), 
	.OE(n2644), 
	.A(\addr_calc/fir_read_addr[11] ));
   TBUFX2TS \addr_calc/addr_tri3[8]  (.Y(addr[8]), 
	.OE(FE_OFN306_n2644), 
	.A(\addr_calc/fir_read_addr[8] ));
   TBUFX2TS \addr_calc/addr_tri3[6]  (.Y(addr[6]), 
	.OE(FE_OFN171_n195), 
	.A(\addr_calc/fir_read_addr[6] ));
   TBUFX2TS \addr_calc/addr_tri3[5]  (.Y(addr[5]), 
	.OE(FE_OFN171_n195), 
	.A(\addr_calc/fir_read_addr[5] ));
   TBUFX16TS \addr_calc/addr_tri4[24]  (.Y(addr[24]), 
	.OE(FE_OFN310_n2643), 
	.A(\addr_calc/fir_write_addr[24] ));
   TBUFX3TS \addr_calc/addr_tri4[20]  (.Y(addr[20]), 
	.OE(FE_OFN173_n131), 
	.A(\addr_calc/fir_write_addr[20] ));
   TBUFX16TS \addr_calc/addr_tri4[17]  (.Y(addr[17]), 
	.OE(FE_OFN172_n131), 
	.A(FE_OFN543_addr_calc_fir_write_addr_17_));
   TBUFX4TS \addr_calc/addr_tri4[14]  (.Y(addr[14]), 
	.OE(n131), 
	.A(\addr_calc/fir_write_addr[14] ));
   TBUFX4TS \addr_calc/addr_tri4[12]  (.Y(addr[12]), 
	.OE(n131), 
	.A(\addr_calc/fir_write_addr[12] ));
   TBUFX3TS \addr_calc/addr_tri4[11]  (.Y(addr[11]), 
	.OE(n2643), 
	.A(\addr_calc/fir_write_addr[11] ));
   TBUFX2TS \addr_calc/addr_tri4[8]  (.Y(addr[8]), 
	.OE(FE_OFN310_n2643), 
	.A(\addr_calc/fir_write_addr[8] ));
   TBUFX2TS \addr_calc/addr_tri4[6]  (.Y(addr[6]), 
	.OE(FE_OFN175_n131), 
	.A(\addr_calc/fir_write_addr[6] ));
   TBUFX2TS \addr_calc/addr_tri4[5]  (.Y(addr[5]), 
	.OE(FE_OFN175_n131), 
	.A(\addr_calc/fir_write_addr[5] ));
   TBUFX16TS \addr_calc/addr_tri5[20]  (.Y(addr[20]), 
	.OE(FE_OFN157_n67), 
	.A(\addr_calc/iir_read_addr[20] ));
   TBUFX8TS \addr_calc/addr_tri5[14]  (.Y(addr[14]), 
	.OE(n67), 
	.A(\addr_calc/iir_read_addr[14] ));
   TBUFX4TS \addr_calc/addr_tri5[12]  (.Y(addr[12]), 
	.OE(n67), 
	.A(\addr_calc/iir_read_addr[12] ));
   TBUFX4TS \addr_calc/addr_tri5[11]  (.Y(addr[11]), 
	.OE(n2642), 
	.A(\addr_calc/iir_read_addr[11] ));
   TBUFX3TS \addr_calc/addr_tri5[8]  (.Y(addr[8]), 
	.OE(FE_OFN294_n2642), 
	.A(\addr_calc/iir_read_addr[8] ));
   TBUFX2TS \addr_calc/addr_tri5[6]  (.Y(addr[6]), 
	.OE(FE_OFN159_n67), 
	.A(\addr_calc/iir_read_addr[6] ));
   TBUFX2TS \addr_calc/addr_tri5[5]  (.Y(addr[5]), 
	.OE(FE_OFN159_n67), 
	.A(\addr_calc/iir_read_addr[5] ));
   TBUFX2TS \addr_calc/addr_tri5[2]  (.Y(addr[2]), 
	.OE(FE_OFN297_n2642), 
	.A(\addr_calc/iir_read_addr[2] ));
   TBUFX4TS \addr_calc/addr_tri6[24]  (.Y(addr[24]), 
	.OE(FE_OFN289_n2641), 
	.A(\addr_calc/iir_write_addr[24] ));
   TBUFX12TS \addr_calc/addr_tri6[20]  (.Y(addr[20]), 
	.OE(FE_OFN153_n3), 
	.A(\addr_calc/iir_write_addr[20] ));
   TBUFX8TS \addr_calc/addr_tri6[17]  (.Y(addr[17]), 
	.OE(FE_OFN152_n3), 
	.A(\addr_calc/iir_write_addr[17] ));
   TBUFX16TS \addr_calc/addr_tri6[14]  (.Y(addr[14]), 
	.OE(n3), 
	.A(\addr_calc/iir_write_addr[14] ));
   TBUFX3TS \addr_calc/addr_tri6[12]  (.Y(addr[12]), 
	.OE(n3), 
	.A(\addr_calc/iir_write_addr[12] ));
   TBUFX3TS \addr_calc/addr_tri6[11]  (.Y(addr[11]), 
	.OE(FE_OFN290_n2641), 
	.A(FE_OFN545_addr_calc_iir_write_addr_11_));
   TBUFX2TS \addr_calc/addr_tri6[8]  (.Y(addr[8]), 
	.OE(FE_OFN290_n2641), 
	.A(\addr_calc/iir_write_addr[8] ));
   TBUFX2TS \addr_calc/addr_tri6[6]  (.Y(addr[6]), 
	.OE(FE_OFN155_n3), 
	.A(\addr_calc/iir_write_addr[6] ));
   TBUFX2TS \addr_calc/addr_tri6[5]  (.Y(addr[5]), 
	.OE(FE_OFN155_n3), 
	.A(\addr_calc/iir_write_addr[5] ));
   DFFQX2TS \addr_calc/fir_read_calc/counter/count_reg[28]  (.Q(\addr_calc/fir_read_calc/count[28] ), 
	.D(n1070), 
	.CK(clk__L1_N0));
   DFFHQX4TS \addr_calc/fir_write_calc/counter/count_reg[2]  (.Q(\addr_calc/fir_write_calc/count[2] ), 
	.D(n1128), 
	.CK(clk__L1_N0));
   DFFX4TS \addr_calc/fir_read_calc/counter/count_reg[29]  (.Q(\addr_calc/fir_read_calc/count[29] ), 
	.D(n1069), 
	.CK(clk__L1_N0));
   DFFHQX2TS \addr_calc/fir_read_calc/counter/count_reg[0]  (.Q(\addr_calc/fir_read_calc/count[0] ), 
	.D(n1098), 
	.CK(clk__L1_N0));
   DFFHQX1TS \addr_calc/iir_read_calc/counter/count_reg[21]  (.Q(\addr_calc/iir_read_calc/count[21] ), 
	.D(n950), 
	.CK(clk__L1_N0));
   DFFHQX1TS \addr_calc/fir_write_calc/counter/count_reg[21]  (.Q(\addr_calc/fir_write_calc/count[21] ), 
	.D(n1109), 
	.CK(clk__L1_N0));
   DFFHQX1TS \addr_calc/fft_write_calc/counter/count_reg[21]  (.Q(\addr_calc/fft_write_calc/count[21] ), 
	.D(n1045), 
	.CK(clk__L1_N0));
   DFFQX1TS \addr_calc/fft_read_calc/counter/count_reg[21]  (.Q(\addr_calc/fft_read_calc/count[21] ), 
	.D(n1013), 
	.CK(clk__L1_N0));
   DFFHQX1TS \addr_calc/fir_write_calc/counter/count_reg[15]  (.Q(\addr_calc/fir_write_calc/count[15] ), 
	.D(n1115), 
	.CK(clk__L1_N0));
   DFFHQX1TS \addr_calc/fir_write_calc/counter/count_reg[19]  (.Q(\addr_calc/fir_write_calc/count[19] ), 
	.D(n1111), 
	.CK(clk__L1_N0));
   DFFHQX2TS \addr_calc/fft_read_calc/counter/count_reg[13]  (.Q(\addr_calc/fft_read_calc/count[13] ), 
	.D(n1021), 
	.CK(clk__L1_N0));
   DFFQX1TS \addr_calc/fft_read_calc/counter/count_reg[17]  (.Q(\addr_calc/fft_read_calc/count[17] ), 
	.D(n1017), 
	.CK(clk__L1_N0));
   DFFHQX2TS \addr_calc/fir_read_calc/counter/count_reg[10]  (.Q(\addr_calc/fir_read_calc/count[10] ), 
	.D(n1088), 
	.CK(clk__L1_N0));
   DFFHQX2TS \addr_calc/fir_read_calc/counter/count_reg[16]  (.Q(\addr_calc/fir_read_calc/count[16] ), 
	.D(n1082), 
	.CK(clk__L1_N0));
   DFFQX1TS \pla_top/fir_enable_reg  (.Q(n2814), 
	.D(n1133), 
	.CK(clk__L1_N0));
   DFFHQX4TS \addr_calc/fft_write_calc/counter/count_reg[4]  (.Q(\addr_calc/fft_write_calc/count[4] ), 
	.D(n1062), 
	.CK(clk__L1_N0));
   DFFHQX2TS \addr_calc/iir_read_calc/counter/count_reg[5]  (.Q(\addr_calc/iir_read_calc/count[5] ), 
	.D(n966), 
	.CK(clk__L1_N0));
   DFFQX4TS \addr_calc/iir_read_calc/counter/count_reg[30]  (.Q(\addr_calc/iir_read_calc/count[30] ), 
	.D(n941), 
	.CK(clk__L1_N0));
   DFFHQX2TS \addr_calc/fir_write_calc/counter/count_reg[14]  (.Q(\addr_calc/fir_write_calc/count[14] ), 
	.D(n1116), 
	.CK(clk__L1_N0));
   DFFHQX2TS \addr_calc/fir_write_calc/counter/count_reg[18]  (.Q(\addr_calc/fir_write_calc/count[18] ), 
	.D(n1112), 
	.CK(clk__L1_N0));
   DFFHQX2TS \addr_calc/fir_read_calc/counter/count_reg[14]  (.Q(\addr_calc/fir_read_calc/count[14] ), 
	.D(n1084), 
	.CK(clk__L1_N0));
   DFFHQX2TS \addr_calc/fir_read_calc/counter/count_reg[18]  (.Q(\addr_calc/fir_read_calc/count[18] ), 
	.D(n1080), 
	.CK(clk__L1_N0));
   DFFHQX2TS \addr_calc/fft_write_calc/counter/count_reg[18]  (.Q(\addr_calc/fft_write_calc/count[18] ), 
	.D(n1048), 
	.CK(clk__L1_N0));
   DFFHQX2TS \addr_calc/fft_read_calc/counter/count_reg[14]  (.Q(\addr_calc/fft_read_calc/count[14] ), 
	.D(n1020), 
	.CK(clk__L1_N0));
   DFFHQX2TS \addr_calc/iir_read_calc/counter/count_reg[18]  (.Q(\addr_calc/iir_read_calc/count[18] ), 
	.D(n953), 
	.CK(clk__L1_N0));
   DFFHQX2TS \addr_calc/fir_write_calc/counter/count_reg[22]  (.Q(\addr_calc/fir_write_calc/count[22] ), 
	.D(n1108), 
	.CK(clk__L1_N0));
   DFFHQX2TS \addr_calc/fir_read_calc/counter/count_reg[22]  (.Q(\addr_calc/fir_read_calc/count[22] ), 
	.D(n1076), 
	.CK(clk__L1_N0));
   DFFQX4TS \addr_calc/fft_write_calc/counter/count_reg[22]  (.Q(\addr_calc/fft_write_calc/count[22] ), 
	.D(n1044), 
	.CK(clk__L1_N0));
   DFFHQX2TS \addr_calc/fft_read_calc/counter/count_reg[22]  (.Q(\addr_calc/fft_read_calc/count[22] ), 
	.D(n1012), 
	.CK(clk__L1_N0));
   DFFQX4TS \addr_calc/fir_write_calc/counter/count_reg[20]  (.Q(\addr_calc/fir_write_calc/count[20] ), 
	.D(n1110), 
	.CK(clk__L1_N0));
   DFFHQX2TS \addr_calc/fir_read_calc/counter/count_reg[20]  (.Q(\addr_calc/fir_read_calc/count[20] ), 
	.D(n1078), 
	.CK(clk__L1_N0));
   DFFQX4TS \addr_calc/fft_write_calc/counter/count_reg[20]  (.Q(\addr_calc/fft_write_calc/count[20] ), 
	.D(n1046), 
	.CK(clk__L1_N0));
   DFFHQX2TS \addr_calc/iir_read_calc/counter/count_reg[20]  (.Q(\addr_calc/iir_read_calc/count[20] ), 
	.D(n951), 
	.CK(clk__L1_N0));
   DFFHQX2TS \addr_calc/fft_read_calc/counter/count_reg[12]  (.Q(\addr_calc/fft_read_calc/count[12] ), 
	.D(n1022), 
	.CK(clk__L1_N0));
   DFFHQX2TS \addr_calc/fft_read_calc/counter/count_reg[0]  (.Q(\addr_calc/fft_read_calc/count[0] ), 
	.D(n1034), 
	.CK(clk__L1_N0));
   DFFHQX4TS \addr_calc/fft_read_calc/counter/count_reg[7]  (.Q(\addr_calc/fft_read_calc/count[7] ), 
	.D(n1027), 
	.CK(clk__L1_N0));
   DFFHQX2TS \addr_calc/iir_write_calc/counter/count_reg[7]  (.Q(\addr_calc/iir_write_calc/count[7] ), 
	.D(n995), 
	.CK(clk__L1_N0));
   DFFHQX2TS \addr_calc/iir_read_calc/counter/count_reg[9]  (.Q(\addr_calc/iir_read_calc/count[9] ), 
	.D(n962), 
	.CK(clk__L1_N0));
   DFFHQX2TS \addr_calc/fir_read_calc/counter/count_reg[30]  (.Q(\addr_calc/fir_read_calc/count[30] ), 
	.D(n1068), 
	.CK(clk__L1_N0));
   DFFX4TS \addr_calc/fft_write_calc/counter/count_reg[30]  (.Q(\addr_calc/fft_write_calc/count[30] ), 
	.D(n1036), 
	.CK(clk__L1_N0));
   DFFHQX8TS \addr_calc/fft_read_calc/counter/count_reg[30]  (.Q(\addr_calc/fft_read_calc/count[30] ), 
	.D(n1004), 
	.CK(clk__L1_N0));
   TBUFX8TS \addr_calc/addr_tri[24]  (.Y(addr[24]), 
	.OE(FE_OFN298_n2646), 
	.A(\addr_calc/fft_read_addr[24] ));
   TBUFX4TS \addr_calc/addr_tri[20]  (.Y(addr[20]), 
	.OE(FE_OFN161_n323), 
	.A(\addr_calc/fft_read_addr[20] ));
   TBUFX16TS \addr_calc/addr_tri[17]  (.Y(addr[17]), 
	.OE(FE_OFN160_n323), 
	.A(\addr_calc/fft_read_addr[17] ));
   AOI21XLTS U346 (.Y(n924), 
	.B0(n925), 
	.A1(n1828), 
	.A0(fir_enable));
   AOI32XLTS U23 (.Y(n791), 
	.B1(FE_OFN228_fft_enable), 
	.B0(fft_read_done), 
	.A2(FE_OFN564_n2066), 
	.A1(FE_OFN561_n2587), 
	.A0(fir_read_done));
   AND2X2TS U342 (.Y(iir_put_req), 
	.B(n796), 
	.A(iir_put_req_reg));
   NOR3XLTS U351 (.Y(n927), 
	.C(n900), 
	.B(n2061), 
	.A(n2071));
   OAI21XLTS U376 (.Y(n939), 
	.B0(n2073), 
	.A1(FE_OFN507_from_fft_empty), 
	.A0(FE_OFN505_to_fft_empty));
   NOR2X2TS U358 (.Y(\data_cntl/N266 ), 
	.B(n2071), 
	.A(FE_OFN565_n2066));
   AOI21X2TS U362 (.Y(\data_cntl/N263 ), 
	.B0(FE_OFN228_fft_enable), 
	.A1(n2061), 
	.A0(iir_enable));
   AOI21XLTS U383 (.Y(n940), 
	.B0(n2072), 
	.A1(FE_OFN563_n2060), 
	.A0(n1861));
   AOI33X1TS U377 (.Y(\data_cntl/N250 ), 
	.B2(FE_OFN506_to_fft_full), 
	.B1(FE_OFN505_to_fft_empty), 
	.B0(n2072), 
	.A2(FE_OFN151_n2074), 
	.A1(FE_OFN507_from_fft_empty), 
	.A0(FE_OFN508_from_fft_full));
   OAI21X1TS U359 (.Y(\data_cntl/N260 ), 
	.B0(FE_OFN561_n2587), 
	.A1(fir_enable), 
	.A0(n2063));
   NOR3X1TS U352 (.Y(n798), 
	.C(n925), 
	.B(FE_OFN563_n2060), 
	.A(n1829));
   NOR3X1TS U25 (.Y(n790), 
	.C(n798), 
	.B(n797), 
	.A(n796));
   AOI31X4TS U21 (.Y(ram_write_enable), 
	.B0(n793), 
	.A2(n792), 
	.A1(n791), 
	.A0(n790));
   NOR2X1TS U314 (.Y(n872), 
	.B(n903), 
	.A(n2311));
   NOR2X1TS U311 (.Y(n902), 
	.B(n903), 
	.A(FE_OFN335_instruction_2_));
   OAI21X1TS U303 (.Y(n873), 
	.B0(n887), 
	.A1(n1828), 
	.A0(fft_read_done));
   AOI21X1TS U301 (.Y(n889), 
	.B0(n884), 
	.A1(n900), 
	.A0(fir_write_done));
   AOI32X1TS U312 (.Y(n891), 
	.B1(FE_OFN146_n801), 
	.B0(n899), 
	.A2(n898), 
	.A1(FE_OFN146_n801), 
	.A0(iir_write_done));
   NOR2X1TS U300 (.Y(n893), 
	.B(n899), 
	.A(n898));
   OAI31X1TS U298 (.Y(n894), 
	.B0(n897), 
	.A2(n1828), 
	.A1(n895), 
	.A0(n870));
   AOI32X1TS U297 (.Y(n892), 
	.B1(FE_OFN146_n801), 
	.B0(n894), 
	.A2(iir_write_done), 
	.A1(n893), 
	.A0(FE_OFN146_n801));
   OAI31X1TS U296 (.Y(n1134), 
	.B0(n892), 
	.A2(n891), 
	.A1(n889), 
	.A0(n890));
   INVX2TS U307 (.Y(n869), 
	.A(FE_OFN145_n801));
   NOR3X1TS U295 (.Y(n886), 
	.C(n889), 
	.B(n888), 
	.A(n887));
   OAI31X1TS U293 (.Y(n1133), 
	.B0(n885), 
	.A2(n884), 
	.A1(n869), 
	.A0(fir_write_done));
   OAI31X1TS U277 (.Y(n1131), 
	.B0(n871), 
	.A2(n870), 
	.A1(n869), 
	.A0(n1478));
   AND2XLTS U379 (.Y(\addr_calc/N223 ), 
	.B(FE_OFN314_data_cntl_N159), 
	.A(\data_cntl/N265 ));
   AND2XLTS U387 (.Y(\addr_calc/N219 ), 
	.B(FE_OFN318_data_cntl_N95), 
	.A(\data_cntl/N262 ));
   AND2XLTS U391 (.Y(\addr_calc/N217 ), 
	.B(FE_OFN322_data_cntl_N9), 
	.A(\data_cntl/N259 ));
   NOR3X1TS U22 (.Y(n793), 
	.C(\data_cntl/N264 ), 
	.B(\data_cntl/N261 ), 
	.A(\data_cntl/N267 ));
   NOR3X1TS U26 (.Y(n795), 
	.C(\data_cntl/N259 ), 
	.B(\data_cntl/N265 ), 
	.A(\data_cntl/N262 ));
   NOR2X4TS U24 (.Y(ram_read_enable), 
	.B(n790), 
	.A(n795));
   NOR2BX1TS U327 (.Y(n801), 
	.B(reset), 
	.AN(chipselect));
   AOI211X4TS U357 (.Y(fft_get_req), 
	.C0(n929), 
	.B0(FE_OFN561_n2587), 
	.A1(n895), 
	.A0(n1829));
   NOR4XLTS U325 (.Y(n904), 
	.D(instruction[25]), 
	.C(instruction[23]), 
	.B(instruction[4]), 
	.A(instruction[5]));
   NOR4XLTS U324 (.Y(n905), 
	.D(instruction[3]), 
	.C(instruction[6]), 
	.B(instruction[7]), 
	.A(instruction[8]));
   NOR4X1TS U339 (.Y(n920), 
	.D(\addr_calc/iir_write_calc/count[20] ), 
	.C(\addr_calc/iir_write_calc/count[21] ), 
	.B(\addr_calc/iir_write_calc/count[22] ), 
	.A(\addr_calc/iir_write_calc/count[23] ));
   NOR4X1TS U337 (.Y(n922), 
	.D(n1945), 
	.C(n2570), 
	.B(FE_OFN230_addr_calc_iir_write_calc_count_15_), 
	.A(n1951));
   NOR4X2TS U72 (.Y(n815), 
	.D(\addr_calc/iir_read_calc/count[20] ), 
	.C(n1687), 
	.B(\addr_calc/iir_read_calc/count[22] ), 
	.A(n2565));
   NOR4X1TS U151 (.Y(n832), 
	.D(FE_OFN287_addr_calc_fft_read_calc_count_17_), 
	.C(\addr_calc/fft_read_calc/count[18] ), 
	.B(\addr_calc/fft_read_calc/count[19] ), 
	.A(n1979));
   NOR4X1TS U150 (.Y(n833), 
	.D(\addr_calc/fft_read_calc/count[20] ), 
	.C(FE_OFN288_addr_calc_fft_read_calc_count_21_), 
	.B(n1665), 
	.A(\addr_calc/fft_read_calc/count[23] ));
   NOR4X2TS U275 (.Y(n866), 
	.D(FE_OFN283_addr_calc_fir_write_calc_count_20_), 
	.C(n1892), 
	.B(n1668), 
	.A(\addr_calc/fir_write_calc/count[23] ));
   NOR4X1TS U273 (.Y(n868), 
	.D(\addr_calc/fir_write_calc/count[13] ), 
	.C(\addr_calc/fir_write_calc/count[14] ), 
	.B(n1883), 
	.A(\addr_calc/fir_write_calc/count[16] ));
   NOR4X2TS U290 (.Y(n881), 
	.D(n1985), 
	.C(n1879), 
	.B(n1691), 
	.A(\addr_calc/fir_read_calc/count[23] ));
   NOR4X1TS U340 (.Y(n919), 
	.D(n1954), 
	.C(FE_OFN266_addr_calc_iir_write_calc_count_18_), 
	.B(\addr_calc/iir_write_calc/count[19] ), 
	.A(n1931));
   NOR4X1TS U73 (.Y(n814), 
	.D(\addr_calc/iir_read_calc/count[17] ), 
	.C(n2025), 
	.B(n2556), 
	.A(n1898));
   NOR4X1TS U196 (.Y(n847), 
	.D(FE_OFN281_addr_calc_fft_write_calc_count_20_), 
	.C(n1918), 
	.B(FE_OFN284_addr_calc_fft_write_calc_count_22_), 
	.A(\addr_calc/fft_write_calc/count[23] ));
   NOR4X1TS U276 (.Y(n865), 
	.D(\addr_calc/fir_write_calc/count[17] ), 
	.C(n2006), 
	.B(\addr_calc/fir_write_calc/count[19] ), 
	.A(\addr_calc/fir_write_calc/count[1] ));
   INVX2TS U353 (.Y(n925), 
	.A(n928));
   DFFHQX8TS \addr_calc/fft_write_calc/counter/count_reg[25]  (.Q(\addr_calc/fft_write_calc/count[25] ), 
	.D(n1041), 
	.CK(clk__L1_N0));
   DFFHQX8TS \addr_calc/iir_write_calc/counter/count_reg[17]  (.Q(\addr_calc/iir_write_calc/count[17] ), 
	.D(n985), 
	.CK(clk__L1_N0));
   DFFHQX8TS \addr_calc/fft_read_calc/counter/count_reg[25]  (.Q(\addr_calc/fft_read_calc/count[25] ), 
	.D(n1009), 
	.CK(clk__L1_N0));
   TBUFX16TS \addr_calc/addr_tri3[30]  (.Y(addr[30]), 
	.OE(FE_OFN308_n2644), 
	.A(\addr_calc/fir_read_addr[30] ));
   DFFHQX8TS \addr_calc/iir_write_calc/counter/count_reg[25]  (.Q(\addr_calc/iir_write_calc/count[25] ), 
	.D(n977), 
	.CK(clk__L1_N0));
   TBUFX16TS \addr_calc/addr_tri5[31]  (.Y(addr[31]), 
	.OE(FE_OFN296_n2642), 
	.A(\addr_calc/iir_read_addr[31] ));
   DFFHQX8TS \addr_calc/fft_read_calc/counter/count_reg[24]  (.Q(\addr_calc/fft_read_calc/count[24] ), 
	.D(n1010), 
	.CK(clk__L1_N0));
   DFFHQX8TS \addr_calc/fir_read_calc/counter/count_reg[25]  (.Q(\addr_calc/fir_read_calc/count[25] ), 
	.D(n1073), 
	.CK(clk__L1_N0));
   DFFHQX4TS \addr_calc/fft_write_calc/counter/count_reg[24]  (.Q(\addr_calc/fft_write_calc/count[24] ), 
	.D(n1042), 
	.CK(clk__L1_N0));
   DFFHQX8TS \addr_calc/iir_read_calc/counter/count_reg[16]  (.Q(\addr_calc/iir_read_calc/count[16] ), 
	.D(n955), 
	.CK(clk__L1_N0));
   TBUFX16TS \addr_calc/addr_tri3[31]  (.Y(addr[31]), 
	.OE(FE_OFN308_n2644), 
	.A(\addr_calc/fir_read_addr[31] ));
   DFFHQX8TS \addr_calc/fir_read_calc/counter/count_reg[24]  (.Q(\addr_calc/fir_read_calc/count[24] ), 
	.D(n1074), 
	.CK(clk__L1_N0));
   DFFHQX8TS \addr_calc/iir_read_calc/counter/count_reg[29]  (.Q(\addr_calc/iir_read_calc/count[29] ), 
	.D(n942), 
	.CK(clk__L1_N0));
   DFFHQX8TS \addr_calc/iir_write_calc/counter/count_reg[19]  (.Q(\addr_calc/iir_write_calc/count[19] ), 
	.D(n983), 
	.CK(clk__L1_N0));
   DFFHQX8TS \addr_calc/iir_read_calc/counter/count_reg[24]  (.Q(\addr_calc/iir_read_calc/count[24] ), 
	.D(n947), 
	.CK(clk__L1_N0));
   TBUFX16TS \addr_calc/addr_tri4[26]  (.Y(addr[26]), 
	.OE(FE_OFN311_n2643), 
	.A(\addr_calc/fir_write_addr[26] ));
   TBUFX12TS \addr_calc/addr_tri4[30]  (.Y(addr[30]), 
	.OE(FE_OFN312_n2643), 
	.A(\addr_calc/fir_write_addr[30] ));
   TBUFX20TS \addr_calc/addr_tri5[27]  (.Y(addr[27]), 
	.OE(FE_OFN295_n2642), 
	.A(\addr_calc/iir_read_addr[27] ));
   DFFHQX8TS \addr_calc/iir_read_calc/counter/count_reg[25]  (.Q(\addr_calc/iir_read_calc/count[25] ), 
	.D(n946), 
	.CK(clk__L1_N0));
   DFFHQX8TS \addr_calc/fft_write_calc/counter/count_reg[29]  (.Q(\addr_calc/fft_write_calc/count[29] ), 
	.D(n1037), 
	.CK(clk__L1_N0));
   DFFHQX4TS \addr_calc/fft_read_calc/counter/count_reg[29]  (.Q(\addr_calc/fft_read_calc/count[29] ), 
	.D(n1005), 
	.CK(clk__L1_N0));
   TBUFX12TS \addr_calc/addr_tri[21]  (.Y(addr[21]), 
	.OE(FE_OFN162_n323), 
	.A(\addr_calc/fft_read_addr[21] ));
   TBUFX16TS \addr_calc/addr_tri4[31]  (.Y(addr[31]), 
	.OE(FE_OFN312_n2643), 
	.A(\addr_calc/fir_write_addr[31] ));
   DFFHQX4TS \addr_calc/iir_write_calc/counter/count_reg[0]  (.Q(\addr_calc/iir_write_calc/count[0] ), 
	.D(n1002), 
	.CK(clk__L1_N0));
   DFFHQX4TS \addr_calc/iir_read_calc/counter/count_reg[3]  (.Q(\addr_calc/iir_read_calc/count[3] ), 
	.D(n968), 
	.CK(clk__L1_N0));
   TBUFX12TS \addr_calc/addr_tri[30]  (.Y(addr[30]), 
	.OE(FE_OFN300_n2646), 
	.A(FE_OFN135_addr_calc_fft_read_addr_30_));
   TBUFX16TS \addr_calc/addr_tri5[30]  (.Y(addr[30]), 
	.OE(FE_OFN296_n2642), 
	.A(\addr_calc/iir_read_addr[30] ));
   DFFHQX4TS \addr_calc/iir_read_calc/counter/count_reg[0]  (.Q(\addr_calc/iir_read_calc/count[0] ), 
	.D(n971), 
	.CK(clk__L1_N0));
   DFFHQX4TS \addr_calc/iir_write_calc/counter/count_reg[5]  (.Q(\addr_calc/iir_write_calc/count[5] ), 
	.D(n997), 
	.CK(clk__L1_N0));
   TBUFX16TS \addr_calc/addr_tri[31]  (.Y(addr[31]), 
	.OE(FE_OFN300_n2646), 
	.A(\addr_calc/fft_read_addr[31] ));
   DFFHQX8TS \addr_calc/fft_read_calc/counter/count_reg[15]  (.Q(\addr_calc/fft_read_calc/count[15] ), 
	.D(n1019), 
	.CK(clk__L1_N0));
   TBUFX12TS \addr_calc/addr_tri6[15]  (.Y(addr[15]), 
	.OE(FE_OFN152_n3), 
	.A(\addr_calc/iir_write_addr[15] ));
   TBUFX16TS \addr_calc/addr_tri4[15]  (.Y(addr[15]), 
	.OE(FE_OFN172_n131), 
	.A(\addr_calc/fir_write_addr[15] ));
   DFFHQX4TS \addr_calc/fft_write_calc/counter/count_reg[31]  (.Q(\addr_calc/fft_write_calc/count[31] ), 
	.D(n1067), 
	.CK(clk__L1_N0));
   DFFHQX4TS \addr_calc/fft_write_calc/counter/count_reg[15]  (.Q(\addr_calc/fft_write_calc/count[15] ), 
	.D(n1051), 
	.CK(clk__L1_N0));
   DFFHQX8TS \addr_calc/fft_write_calc/counter/count_reg[27]  (.Q(\addr_calc/fft_write_calc/count[27] ), 
	.D(n1039), 
	.CK(clk__L1_N0));
   TBUFX16TS \addr_calc/addr_tri4[23]  (.Y(addr[23]), 
	.OE(FE_OFN174_n131), 
	.A(\addr_calc/fir_write_addr[23] ));
   DFFHQX4TS \addr_calc/fft_read_calc/counter/count_reg[19]  (.Q(\addr_calc/fft_read_calc/count[19] ), 
	.D(n1015), 
	.CK(clk__L1_N0));
   TBUFX16TS \addr_calc/addr_tri[26]  (.Y(addr[26]), 
	.OE(FE_OFN299_n2646), 
	.A(\addr_calc/fft_read_addr[26] ));
   TBUFX16TS \addr_calc/addr_tri5[26]  (.Y(addr[26]), 
	.OE(FE_OFN295_n2642), 
	.A(\addr_calc/iir_read_addr[26] ));
   TBUFX12TS \addr_calc/addr_tri6[26]  (.Y(addr[26]), 
	.OE(FE_OFN291_n2641), 
	.A(\addr_calc/iir_write_addr[26] ));
   TBUFX8TS \addr_calc/addr_tri3[26]  (.Y(addr[26]), 
	.OE(FE_OFN307_n2644), 
	.A(\addr_calc/fir_read_addr[26] ));
   DFFHQX4TS \addr_calc/fir_write_calc/counter/count_reg[9]  (.Q(\addr_calc/fir_write_calc/count[9] ), 
	.D(n1121), 
	.CK(clk__L1_N0));
   TBUFX8TS \addr_calc/addr_tri4[22]  (.Y(addr[22]), 
	.OE(FE_OFN174_n131), 
	.A(\addr_calc/fir_write_addr[22] ));
   DFFHQX4TS \addr_calc/iir_write_calc/counter/count_reg[27]  (.Q(\addr_calc/iir_write_calc/count[27] ), 
	.D(n975), 
	.CK(clk__L1_N0));
   DFFHQX8TS \addr_calc/fir_write_calc/counter/count_reg[29]  (.Q(\addr_calc/fir_write_calc/count[29] ), 
	.D(n1101), 
	.CK(clk__L1_N0));
   DFFHQX8TS \addr_calc/fft_write_calc/counter/count_reg[6]  (.Q(\addr_calc/fft_write_calc/count[6] ), 
	.D(n1060), 
	.CK(clk__L1_N0));
   DFFHQX4TS \addr_calc/fft_write_calc/counter/count_reg[13]  (.Q(\addr_calc/fft_write_calc/count[13] ), 
	.D(n1053), 
	.CK(clk__L1_N0));
   DFFHQX4TS \addr_calc/iir_write_calc/counter/count_reg[21]  (.Q(\addr_calc/iir_write_calc/count[21] ), 
	.D(n981), 
	.CK(clk__L1_N0));
   DFFHQX4TS \addr_calc/iir_write_calc/counter/count_reg[28]  (.Q(\addr_calc/iir_write_calc/count[28] ), 
	.D(n974), 
	.CK(clk__L1_N0));
   DFFHQX2TS \addr_calc/fir_write_calc/counter/count_reg[27]  (.Q(\addr_calc/fir_write_calc/count[27] ), 
	.D(n1103), 
	.CK(clk__L1_N0));
   DFFHQX4TS \addr_calc/fir_write_calc/counter/count_reg[17]  (.Q(\addr_calc/fir_write_calc/count[17] ), 
	.D(n1113), 
	.CK(clk__L1_N0));
   DFFHQX4TS \addr_calc/fir_write_calc/counter/count_reg[5]  (.Q(\addr_calc/fir_write_calc/count[5] ), 
	.D(n1125), 
	.CK(clk__L1_N0));
   DFFHQX4TS \addr_calc/fft_write_calc/counter/count_reg[11]  (.Q(\addr_calc/fft_write_calc/count[11] ), 
	.D(n1055), 
	.CK(clk__L1_N0));
   DFFHQX4TS \addr_calc/fft_read_calc/counter/count_reg[27]  (.Q(\addr_calc/fft_read_calc/count[27] ), 
	.D(n1007), 
	.CK(clk__L1_N0));
   DFFHQX4TS \addr_calc/fft_write_calc/counter/count_reg[19]  (.Q(\addr_calc/fft_write_calc/count[19] ), 
	.D(n1047), 
	.CK(clk__L1_N0));
   OAI21X1TS \add_x_19_4/U70  (.Y(\add_x_19_4/n77 ), 
	.B0(\add_x_19_4/n79 ), 
	.A1(\add_x_19_4/n82 ), 
	.A0(\add_x_19_4/n78 ));
   NAND2X2TS \add_x_19_4/U255  (.Y(\add_x_19_4/n191 ), 
	.B(FE_OCPUNCON1077_FE_OFN459_offset_0_), 
	.A(\addr_calc/iir_read_calc/count[0] ));
   XOR2X1TS \add_x_19_4/U244  (.Y(\addr_calc/iir_read_addr[1] ), 
	.B(\add_x_19_4/n191 ), 
	.A(\add_x_19_4/n31 ));
   XOR2X1TS \add_x_19_4/U238  (.Y(\addr_calc/iir_read_addr[2] ), 
	.B(\add_x_19_4/n30 ), 
	.A(\add_x_19_4/n186 ));
   AOI21X2TS \add_x_19_4/U214  (.Y(\add_x_19_4/n167 ), 
	.B0(\add_x_19_4/n169 ), 
	.A1(\add_x_19_4/n168 ), 
	.A0(FE_OCP_RBN1978_add_x_19_4_n178));
   AOI21X4TS \add_x_19_4/U173  (.Y(\add_x_19_4/n141 ), 
	.B0(\add_x_19_4/n143 ), 
	.A1(\add_x_19_4/n213 ), 
	.A0(\add_x_19_4/n146 ));
   OAI21X4TS \add_x_19_4/U156  (.Y(\add_x_19_4/n130 ), 
	.B0(\add_x_19_4/n132 ), 
	.A1(\add_x_19_4/n131 ), 
	.A0(\add_x_19_4/n133 ));
   OAI21X2TS \add_x_19_4/U90  (.Y(\add_x_19_4/n88 ), 
	.B0(\add_x_19_4/n90 ), 
	.A1(\add_x_19_4/n89 ), 
	.A0(\add_x_19_4/n91 ));
   NOR2X1TS \add_x_19_4/U10  (.Y(\add_x_19_4/n36 ), 
	.B(FE_OFN559_offset_30_), 
	.A(FE_OFN286_addr_calc_iir_read_calc_count_30_));
   AOI21X2TS \add_x_19_4/U33  (.Y(\add_x_19_4/n52 ), 
	.B0(\add_x_19_4/n54 ), 
	.A1(\add_x_19_4/n62 ), 
	.A0(\add_x_19_4/n53 ));
   OAI21X2TS \add_x_19_4/U35  (.Y(\add_x_19_4/n54 ), 
	.B0(\add_x_19_4/n56 ), 
	.A1(\add_x_19_4/n59 ), 
	.A0(\add_x_19_4/n55 ));
   OAI21X2TS \add_x_19_4/U49  (.Y(\add_x_19_4/n62 ), 
	.B0(\add_x_19_4/n64 ), 
	.A1(\add_x_19_4/n67 ), 
	.A0(\add_x_19_4/n63 ));
   OAI21X2TS \add_x_19_4/U84  (.Y(\add_x_19_4/n85 ), 
	.B0(\add_x_19_4/n87 ), 
	.A1(\add_x_19_4/n90 ), 
	.A0(\add_x_19_4/n86 ));
   AOI21X4TS \add_x_19_4/U99  (.Y(\add_x_19_4/n94 ), 
	.B0(\add_x_19_4/n96 ), 
	.A1(\add_x_19_4/n104 ), 
	.A0(\add_x_19_4/n95 ));
   OAI21X2TS \add_x_19_4/U101  (.Y(\add_x_19_4/n96 ), 
	.B0(\add_x_19_4/n98 ), 
	.A1(\add_x_19_4/n101 ), 
	.A0(\add_x_19_4/n97 ));
   NOR2X2TS \add_x_19_4/U24  (.Y(\add_x_19_4/n46 ), 
	.B(\add_x_19_4/n48 ), 
	.A(\add_x_19_4/n51 ));
   NOR2X1TS \add_x_19_4/U34  (.Y(\add_x_19_4/n53 ), 
	.B(\add_x_19_4/n55 ), 
	.A(\add_x_19_4/n58 ));
   NOR2X1TS \add_x_19_4/U83  (.Y(\add_x_19_4/n84 ), 
	.B(\add_x_19_4/n89 ), 
	.A(\add_x_19_4/n86 ));
   NOR2X1TS \add_x_19_4/U100  (.Y(\add_x_19_4/n95 ), 
	.B(\add_x_19_4/n97 ), 
	.A(\add_x_19_4/n100 ));
   NOR2X4TS \add_x_19_4/U114  (.Y(\add_x_19_4/n103 ), 
	.B(\add_x_19_4/n105 ), 
	.A(\add_x_19_4/n110 ));
   OAI21X2TS \add_x_19_4/U167  (.Y(\add_x_19_4/n138 ), 
	.B0(\add_x_19_4/n140 ), 
	.A1(\add_x_19_4/n145 ), 
	.A0(\add_x_19_4/n139 ));
   NOR2X2TS \add_x_19_4/U166  (.Y(\add_x_19_4/n137 ), 
	.B(\add_x_19_4/n139 ), 
	.A(\add_x_19_4/n144 ));
   NOR2X1TS \add_x_19_4/U184  (.Y(\add_x_19_4/n149 ), 
	.B(\add_x_19_4/n151 ), 
	.A(\add_x_19_4/n154 ));
   NOR2X8TS \add_x_19_4/U201  (.Y(\add_x_19_4/n160 ), 
	.B(\add_x_19_4/n162 ), 
	.A(\add_x_19_4/n165 ));
   NOR2X4TS \add_x_19_4/U215  (.Y(\add_x_19_4/n168 ), 
	.B(\add_x_19_4/n170 ), 
	.A(\add_x_19_4/n175 ));
   NOR2X2TS \add_x_19_4/U249  (.Y(\add_x_19_4/n188 ), 
	.B(FE_OCP_RBN1919_offset_1_), 
	.A(\addr_calc/iir_read_calc/count[1] ));
   XOR2X2TS \add_x_19_4/U207  (.Y(\addr_calc/iir_read_addr[6] ), 
	.B(\add_x_19_4/n26 ), 
	.A(\add_x_19_4/n167 ));
   XOR2X4TS \add_x_19_4/U161  (.Y(\addr_calc/iir_read_addr[11] ), 
	.B(\add_x_19_4/n21 ), 
	.A(\add_x_19_4/n141 ));
   NAND2X1TS \add_x_19_4/U11  (.Y(\add_x_19_4/n37 ), 
	.B(FE_OFN559_offset_30_), 
	.A(FE_OFN286_addr_calc_iir_read_calc_count_30_));
   NAND2X1TS \add_x_19_4/U19  (.Y(\add_x_19_4/n42 ), 
	.B(FE_OFN347_offset_29_), 
	.A(n1840));
   NAND2X1TS \add_x_19_4/U29  (.Y(\add_x_19_4/n49 ), 
	.B(FE_OFN351_offset_28_), 
	.A(n2561));
   NAND2X1TS \add_x_19_4/U39  (.Y(\add_x_19_4/n56 ), 
	.B(FE_OFN355_offset_27_), 
	.A(FE_OFN235_addr_calc_iir_read_calc_count_27_));
   NAND2X1TS \add_x_19_4/U45  (.Y(\add_x_19_4/n59 ), 
	.B(FE_OFN360_offset_26_), 
	.A(\addr_calc/iir_read_calc/count[26] ));
   NAND2X1TS \add_x_19_4/U53  (.Y(\add_x_19_4/n64 ), 
	.B(FE_OFN364_offset_25_), 
	.A(n1926));
   NAND2X1TS \add_x_19_4/U59  (.Y(\add_x_19_4/n67 ), 
	.B(FE_OFN367_offset_24_), 
	.A(n2034));
   NAND2X1TS \add_x_19_4/U74  (.Y(\add_x_19_4/n79 ), 
	.B(FE_OFN372_offset_23_), 
	.A(\addr_calc/iir_read_calc/count[23] ));
   NAND2X1TS \add_x_19_4/U80  (.Y(\add_x_19_4/n82 ), 
	.B(FE_OCPUNCON1877_FE_OFN374_offset_22_), 
	.A(\addr_calc/iir_read_calc/count[22] ));
   NAND2X1TS \add_x_19_4/U88  (.Y(\add_x_19_4/n87 ), 
	.B(FE_OFN380_offset_21_), 
	.A(n1687));
   NAND2X1TS \add_x_19_4/U94  (.Y(\add_x_19_4/n90 ), 
	.B(FE_OFN558_n2441), 
	.A(n2028));
   NAND2X1TS \add_x_19_4/U105  (.Y(\add_x_19_4/n98 ), 
	.B(FE_OFN384_offset_19_), 
	.A(\addr_calc/iir_read_calc/count[19] ));
   NAND2X1TS \add_x_19_4/U111  (.Y(\add_x_19_4/n101 ), 
	.B(FE_OFN389_offset_18_), 
	.A(n2025));
   NAND2X6TS \add_x_19_4/U127  (.Y(\add_x_19_4/n111 ), 
	.B(FE_OFN397_offset_16_), 
	.A(n1916));
   NOR2X2TS \add_x_19_4/U58  (.Y(\add_x_19_4/n66 ), 
	.B(FE_OFN367_offset_24_), 
	.A(\addr_calc/iir_read_calc/count[24] ));
   NOR2X6TS \add_x_19_4/U87  (.Y(\add_x_19_4/n86 ), 
	.B(n1687), 
	.A(FE_OFN380_offset_21_));
   NOR2X6TS \add_x_19_4/U93  (.Y(\add_x_19_4/n89 ), 
	.B(n2028), 
	.A(FE_OFN558_n2441));
   NOR2X4TS \add_x_19_4/U110  (.Y(\add_x_19_4/n100 ), 
	.B(FE_OFN389_offset_18_), 
	.A(n2025));
   NOR2X6TS \add_x_19_4/U118  (.Y(\add_x_19_4/n105 ), 
	.B(FE_OFN392_offset_17_), 
	.A(n1920));
   NOR2X1TS \add_x_19_4/U126  (.Y(\add_x_19_4/n110 ), 
	.B(FE_OFN397_offset_16_), 
	.A(n1916));
   NAND2X1TS \add_x_19_4/U140  (.Y(\add_x_19_4/n121 ), 
	.B(FE_OCPUNCON1942_FE_OFN399_offset_15_), 
	.A(\addr_calc/iir_read_calc/count[15] ));
   NAND2X1TS \add_x_19_4/U154  (.Y(\add_x_19_4/n129 ), 
	.B(FE_OFN408_offset_13_), 
	.A(\addr_calc/iir_read_calc/count[13] ));
   NAND2X1TS \add_x_19_4/U179  (.Y(\add_x_19_4/n145 ), 
	.B(FE_OFN421_offset_10_), 
	.A(FE_OFN248_addr_calc_iir_read_calc_count_10_));
   NAND2X1TS \add_x_19_4/U189  (.Y(\add_x_19_4/n152 ), 
	.B(FE_OFN424_offset_9_), 
	.A(n1685));
   NAND2X1TS \add_x_19_4/U195  (.Y(\add_x_19_4/n155 ), 
	.B(FE_OFN429_offset_8_), 
	.A(\addr_calc/iir_read_calc/count[8] ));
   NOR2X2TS \add_x_19_4/U153  (.Y(\add_x_19_4/n128 ), 
	.B(FE_OFN408_offset_13_), 
	.A(\addr_calc/iir_read_calc/count[13] ));
   NOR2X1TS \add_x_19_4/U178  (.Y(\add_x_19_4/n144 ), 
	.B(FE_OFN421_offset_10_), 
	.A(FE_OFN248_addr_calc_iir_read_calc_count_10_));
   NOR2X1TS \add_x_19_4/U194  (.Y(\add_x_19_4/n154 ), 
	.B(FE_OFN429_offset_8_), 
	.A(\addr_calc/iir_read_calc/count[8] ));
   NAND2X4TS \add_x_19_4/U206  (.Y(\add_x_19_4/n163 ), 
	.B(FE_OCP_RBN1840_offset_7_), 
	.A(FE_OFN247_addr_calc_iir_read_calc_count_7_));
   NAND2X1TS \add_x_19_4/U212  (.Y(\add_x_19_4/n166 ), 
	.B(\addr_calc/iir_read_calc/count[6] ), 
	.A(FE_OFN436_offset_6_));
   NAND2X2TS \add_x_19_4/U228  (.Y(\add_x_19_4/n176 ), 
	.B(FE_OFN444_offset_4_), 
	.A(FE_OFN244_addr_calc_iir_read_calc_count_4_));
   NOR2X2TS \add_x_19_4/U211  (.Y(\add_x_19_4/n165 ), 
	.B(FE_OFN436_offset_6_), 
	.A(\addr_calc/iir_read_calc/count[6] ));
   NOR2X2TS \add_x_19_4/U227  (.Y(\add_x_19_4/n175 ), 
	.B(FE_OFN444_offset_4_), 
	.A(FE_OFN244_addr_calc_iir_read_calc_count_4_));
   NAND2X1TS \add_x_19_4/U237  (.Y(\add_x_19_4/n182 ), 
	.B(FE_OCPUNCON1075_FE_OFN447_offset_3_), 
	.A(n1902));
   NAND2X1TS \add_x_19_4/U250  (.Y(\add_x_19_4/n189 ), 
	.B(\addr_calc/iir_read_calc/count[1] ), 
	.A(FE_OCP_RBN1919_offset_1_));
   NOR2X2TS \add_x_19_4/U242  (.Y(\add_x_19_4/n184 ), 
	.B(FE_OCPUNCON1076_FE_OFN451_offset_2_), 
	.A(\addr_calc/iir_read_calc/count[2] ));
   NAND2X1TS \add_x_19_4/U247  (.Y(\add_x_19_4/n31 ), 
	.B(\add_x_19_4/n189 ), 
	.A(\add_x_19_4/n222 ));
   NAND2X1TS \add_x_19_4/U240  (.Y(\add_x_19_4/n30 ), 
	.B(\add_x_19_4/n185 ), 
	.A(\add_x_19_4/n221 ));
   XNOR2XLTS \add_x_19_4/U221  (.Y(\addr_calc/iir_read_addr[4] ), 
	.B(\add_x_19_4/n28 ), 
	.A(FE_OCP_RBN1978_add_x_19_4_n178));
   NAND2X1TS \add_x_19_4/U225  (.Y(\add_x_19_4/n28 ), 
	.B(\add_x_19_4/n176 ), 
	.A(\add_x_19_4/n219 ));
   NAND2X1TS \add_x_19_4/U209  (.Y(\add_x_19_4/n26 ), 
	.B(\add_x_19_4/n166 ), 
	.A(\add_x_19_4/n217 ));
   XNOR2X1TS \add_x_19_4/U172  (.Y(\addr_calc/iir_read_addr[10] ), 
	.B(\add_x_19_4/n22 ), 
	.A(\add_x_19_4/n146 ));
   NAND2X1TS \add_x_19_4/U176  (.Y(\add_x_19_4/n22 ), 
	.B(\add_x_19_4/n145 ), 
	.A(\add_x_19_4/n213 ));
   NAND2X1TS \add_x_19_4/U168  (.Y(\add_x_19_4/n21 ), 
	.B(\add_x_19_4/n140 ), 
	.A(\add_x_19_4/n212 ));
   XNOR2X4TS \add_x_19_4/U147  (.Y(\addr_calc/iir_read_addr[13] ), 
	.B(\add_x_19_4/n19 ), 
	.A(\add_x_19_4/n130 ));
   NAND2X1TS \add_x_19_4/U151  (.Y(\add_x_19_4/n19 ), 
	.B(\add_x_19_4/n129 ), 
	.A(n1632));
   NAND2X1TS \add_x_19_4/U116  (.Y(\add_x_19_4/n15 ), 
	.B(\add_x_19_4/n106 ), 
	.A(\add_x_19_4/n206 ));
   XNOR2X4TS \add_x_19_4/U12  (.Y(\addr_calc/iir_read_addr[29] ), 
	.B(\add_x_19_4/n3 ), 
	.A(FE_OCPUNCON1650_add_x_19_4_n43));
   NAND2X1TS \add_x_19_4/U16  (.Y(\add_x_19_4/n3 ), 
	.B(\add_x_19_4/n42 ), 
	.A(n2634));
   NAND2X1TS \add_x_19_4/U102  (.Y(\add_x_19_4/n13 ), 
	.B(\add_x_19_4/n98 ), 
	.A(\add_x_19_4/n204 ));
   NAND2XLTS \add_x_19_4/U85  (.Y(\add_x_19_4/n11 ), 
	.B(\add_x_19_4/n87 ), 
	.A(\add_x_19_4/n202 ));
   NAND2X1TS \add_x_19_4/U36  (.Y(\add_x_19_4/n5 ), 
	.B(\add_x_19_4/n56 ), 
	.A(\add_x_19_4/n196 ));
   NAND2X1TS \add_x_19_4/U119  (.Y(\add_x_19_4/n106 ), 
	.B(FE_OFN392_offset_17_), 
	.A(n1920));
   NAND2X1TS \add_x_19_4/U32  (.Y(\add_x_19_4/n51 ), 
	.B(\add_x_19_4/n53 ), 
	.A(\add_x_19_4/n61 ));
   NAND2X4TS \add_x_19_4/U98  (.Y(\add_x_19_4/n93 ), 
	.B(\add_x_19_4/n95 ), 
	.A(\add_x_19_4/n103 ));
   NAND2X1TS \add_x_19_4/U171  (.Y(\add_x_19_4/n140 ), 
	.B(FE_OFN417_offset_11_), 
	.A(FE_OFN237_addr_calc_iir_read_calc_count_11_));
   NAND2X2TS \add_x_19_4/U164  (.Y(\add_x_19_4/n135 ), 
	.B(\add_x_19_4/n137 ), 
	.A(\add_x_19_4/n149 ));
   NAND2X2TS \add_x_19_4/U220  (.Y(\add_x_19_4/n171 ), 
	.B(FE_OCP_RBN1492_offset_5_), 
	.A(\addr_calc/iir_read_calc/count[5] ));
   NOR2X8TS \add_x_19_2/U236  (.Y(\add_x_19_2/n181 ), 
	.B(FE_OCPN1904_FE_OCPUNCON1066_offset_3_), 
	.A(\addr_calc/fir_read_calc/count[3] ));
   NOR2X6TS \add_x_19_2/U211  (.Y(\add_x_19_2/n165 ), 
	.B(FE_OFN435_offset_6_), 
	.A(\addr_calc/fir_read_calc/count[6] ));
   NAND2X6TS \add_x_19_2/U255  (.Y(\add_x_19_2/n191 ), 
	.B(\addr_calc/fir_read_calc/count[0] ), 
	.A(FE_OCPUNCON1068_offset_0_));
   OAI21X1TS \add_x_19_2/U208  (.Y(\add_x_19_2/n164 ), 
	.B0(\add_x_19_2/n166 ), 
	.A1(\add_x_19_2/n165 ), 
	.A0(\add_x_19_2/n167 ));
   AOI21X1TS \add_x_19_2/U214  (.Y(\add_x_19_2/n167 ), 
	.B0(\add_x_19_2/n169 ), 
	.A1(\add_x_19_2/n168 ), 
	.A0(\add_x_19_2/n177 ));
   OAI21X2TS \add_x_19_2/U181  (.Y(\add_x_19_2/n146 ), 
	.B0(\add_x_19_2/n148 ), 
	.A1(\add_x_19_2/n147 ), 
	.A0(\add_x_19_2/n156 ));
   AOI21X4TS \add_x_19_2/U121  (.Y(\add_x_19_2/n107 ), 
	.B0(\add_x_19_2/n109 ), 
	.A1(\add_x_19_2/n207 ), 
	.A0(\add_x_19_2/n112 ));
   OAI21X1TS \add_x_19_2/U142  (.Y(\add_x_19_2/n122 ), 
	.B0(\add_x_19_2/n124 ), 
	.A1(\add_x_19_2/n123 ), 
	.A0(\add_x_19_2/n125 ));
   AOI21X4TS \add_x_19_2/U148  (.Y(\add_x_19_2/n125 ), 
	.B0(\add_x_19_2/n127 ), 
	.A1(\add_x_19_2/n134 ), 
	.A0(\add_x_19_2/n126 ));
   AOI21X2TS \add_x_19_2/U113  (.Y(\add_x_19_2/n102 ), 
	.B0(\add_x_19_2/n104 ), 
	.A1(\add_x_19_2/n103 ), 
	.A0(\add_x_19_2/n112 ));
   NOR2X1TS \add_x_19_2/U10  (.Y(\add_x_19_2/n36 ), 
	.B(FE_OFN343_offset_30_), 
	.A(n1838));
   OAI21X2TS \add_x_19_2/U49  (.Y(\add_x_19_2/n62 ), 
	.B0(\add_x_19_2/n64 ), 
	.A1(\add_x_19_2/n67 ), 
	.A0(\add_x_19_2/n63 ));
   OAI21X1TS \add_x_19_2/U101  (.Y(\add_x_19_2/n96 ), 
	.B0(\add_x_19_2/n98 ), 
	.A1(\add_x_19_2/n101 ), 
	.A0(\add_x_19_2/n97 ));
   NOR2X1TS \add_x_19_2/U48  (.Y(\add_x_19_2/n61 ), 
	.B(\add_x_19_2/n63 ), 
	.A(\add_x_19_2/n66 ));
   NOR2X1TS \add_x_19_2/U58  (.Y(\add_x_19_2/n66 ), 
	.B(FE_OFN366_offset_24_), 
	.A(n1983));
   NOR2X4TS \add_x_19_2/U65  (.Y(\add_x_19_2/n72 ), 
	.B(\add_x_19_2/n74 ), 
	.A(\add_x_19_2/n93 ));
   NOR2X2TS \add_x_19_2/U83  (.Y(\add_x_19_2/n84 ), 
	.B(\add_x_19_2/n86 ), 
	.A(\add_x_19_2/n89 ));
   NOR2X1TS \add_x_19_2/U100  (.Y(\add_x_19_2/n95 ), 
	.B(\add_x_19_2/n97 ), 
	.A(\add_x_19_2/n100 ));
   NOR2X1TS \add_x_19_2/U114  (.Y(\add_x_19_2/n103 ), 
	.B(\add_x_19_2/n105 ), 
	.A(\add_x_19_2/n110 ));
   OAI21X2TS \add_x_19_2/U150  (.Y(\add_x_19_2/n127 ), 
	.B0(\add_x_19_2/n129 ), 
	.A1(\add_x_19_2/n132 ), 
	.A0(\add_x_19_2/n128 ));
   NOR2X1TS \add_x_19_2/U139  (.Y(\add_x_19_2/n120 ), 
	.B(FE_OCPUNCON1940_offset_15_), 
	.A(\addr_calc/fir_read_calc/count[15] ));
   NOR2X2TS \add_x_19_2/U149  (.Y(\add_x_19_2/n126 ), 
	.B(\add_x_19_2/n128 ), 
	.A(\add_x_19_2/n131 ));
   NOR2X2TS \add_x_19_2/U166  (.Y(\add_x_19_2/n137 ), 
	.B(\add_x_19_2/n139 ), 
	.A(\add_x_19_2/n144 ));
   NOR2X1TS \add_x_19_2/U170  (.Y(\add_x_19_2/n139 ), 
	.B(FE_OCPUNCON652_FE_OFN414_offset_11_), 
	.A(\addr_calc/fir_read_calc/count[11] ));
   NOR2X1TS \add_x_19_2/U184  (.Y(\add_x_19_2/n149 ), 
	.B(\add_x_19_2/n151 ), 
	.A(\add_x_19_2/n154 ));
   NOR2X2TS \add_x_19_2/U215  (.Y(\add_x_19_2/n168 ), 
	.B(\add_x_19_2/n175 ), 
	.A(\add_x_19_2/n170 ));
   NOR2X1TS \add_x_19_2/U249  (.Y(\add_x_19_2/n188 ), 
	.B(FE_OFN249_addr_calc_fir_read_calc_count_1_), 
	.A(FE_OCP_RBN1974_offset_1_));
   NAND2X1TS \add_x_19_2/U11  (.Y(\add_x_19_2/n37 ), 
	.B(FE_OFN343_offset_30_), 
	.A(\addr_calc/fir_read_calc/count[30] ));
   NAND2X1TS \add_x_19_2/U19  (.Y(\add_x_19_2/n42 ), 
	.B(FE_OFN346_offset_29_), 
	.A(n1842));
   NAND2X1TS \add_x_19_2/U29  (.Y(\add_x_19_2/n49 ), 
	.B(FE_OFN350_offset_28_), 
	.A(n1871));
   NAND2X1TS \add_x_19_2/U39  (.Y(\add_x_19_2/n56 ), 
	.B(FE_OFN354_offset_27_), 
	.A(\addr_calc/fir_read_calc/count[27] ));
   NAND2X1TS \add_x_19_2/U45  (.Y(\add_x_19_2/n59 ), 
	.B(FE_OFN357_offset_26_), 
	.A(FE_OFN269_addr_calc_fir_read_calc_count_26_));
   NAND2X1TS \add_x_19_2/U53  (.Y(\add_x_19_2/n64 ), 
	.B(FE_OCPUNCON1318_FE_OFN361_offset_25_), 
	.A(n1876));
   NAND2X1TS \add_x_19_2/U59  (.Y(\add_x_19_2/n67 ), 
	.B(FE_OFN366_offset_24_), 
	.A(n1983));
   NAND2X1TS \add_x_19_2/U74  (.Y(\add_x_19_2/n79 ), 
	.B(FE_OFN369_offset_23_), 
	.A(\addr_calc/fir_read_calc/count[23] ));
   NAND2X1TS \add_x_19_2/U80  (.Y(\add_x_19_2/n82 ), 
	.B(FE_OCPUNCON1876_offset_22_), 
	.A(\addr_calc/fir_read_calc/count[22] ));
   NAND2X1TS \add_x_19_2/U88  (.Y(\add_x_19_2/n87 ), 
	.B(FE_OCPUNCON1070_FE_OFN377_offset_21_), 
	.A(n1879));
   NAND2X1TS \add_x_19_2/U94  (.Y(\add_x_19_2/n90 ), 
	.B(n2441), 
	.A(n1985));
   NAND2X1TS \add_x_19_2/U105  (.Y(\add_x_19_2/n98 ), 
	.B(FE_OCPUNCON1071_FE_OFN382_offset_19_), 
	.A(\addr_calc/fir_read_calc/count[19] ));
   NAND2X1TS \add_x_19_2/U111  (.Y(\add_x_19_2/n101 ), 
	.B(FE_OCPUNCON1072_FE_OFN386_offset_18_), 
	.A(n1988));
   NAND2X1TS \add_x_19_2/U127  (.Y(\add_x_19_2/n111 ), 
	.B(FE_OFN394_offset_16_), 
	.A(n1888));
   NOR2X1TS \add_x_19_2/U52  (.Y(\add_x_19_2/n63 ), 
	.B(FE_OCPUNCON1318_FE_OFN361_offset_25_), 
	.A(n1876));
   NOR2X1TS \add_x_19_2/U79  (.Y(\add_x_19_2/n81 ), 
	.B(FE_OCPUNCON1876_offset_22_), 
	.A(n1691));
   NOR2X1TS \add_x_19_2/U93  (.Y(\add_x_19_2/n89 ), 
	.B(n1985), 
	.A(FE_OFN557_n2441));
   NOR2X1TS \add_x_19_2/U104  (.Y(\add_x_19_2/n97 ), 
	.B(FE_OCPUNCON1071_FE_OFN382_offset_19_), 
	.A(\addr_calc/fir_read_calc/count[19] ));
   NOR2X1TS \add_x_19_2/U110  (.Y(\add_x_19_2/n100 ), 
	.B(FE_OCPUNCON1072_FE_OFN386_offset_18_), 
	.A(n1988));
   NOR2X6TS \add_x_19_2/U118  (.Y(\add_x_19_2/n105 ), 
	.B(FE_OFN391_offset_17_), 
	.A(\addr_calc/fir_read_calc/count[17] ));
   NOR2X1TS \add_x_19_2/U126  (.Y(\add_x_19_2/n110 ), 
	.B(FE_OFN394_offset_16_), 
	.A(n1888));
   NAND2X1TS \add_x_19_2/U140  (.Y(\add_x_19_2/n121 ), 
	.B(FE_OCPUNCON1940_offset_15_), 
	.A(\addr_calc/fir_read_calc/count[15] ));
   NAND2X1TS \add_x_19_2/U146  (.Y(\add_x_19_2/n124 ), 
	.B(FE_OFN402_offset_14_), 
	.A(\addr_calc/fir_read_calc/count[14] ));
   NAND2X1TS \add_x_19_2/U154  (.Y(\add_x_19_2/n129 ), 
	.B(FE_OFN407_offset_13_), 
	.A(\addr_calc/fir_read_calc/count[13] ));
   NAND2X1TS \add_x_19_2/U160  (.Y(\add_x_19_2/n132 ), 
	.B(FE_OFN411_offset_12_), 
	.A(\addr_calc/fir_read_calc/count[12] ));
   NAND2X1TS \add_x_19_2/U189  (.Y(\add_x_19_2/n152 ), 
	.B(FE_OCPUNCON654_FE_OFN422_offset_9_), 
	.A(n1900));
   NAND2X1TS \add_x_19_2/U195  (.Y(\add_x_19_2/n155 ), 
	.B(FE_OFN426_offset_8_), 
	.A(\addr_calc/fir_read_calc/count[8] ));
   NOR2X1TS \add_x_19_2/U153  (.Y(\add_x_19_2/n128 ), 
	.B(FE_OFN407_offset_13_), 
	.A(\addr_calc/fir_read_calc/count[13] ));
   NOR2X1TS \add_x_19_2/U159  (.Y(\add_x_19_2/n131 ), 
	.B(FE_OFN411_offset_12_), 
	.A(\addr_calc/fir_read_calc/count[12] ));
   NOR2X1TS \add_x_19_2/U194  (.Y(\add_x_19_2/n154 ), 
	.B(FE_OFN426_offset_8_), 
	.A(\addr_calc/fir_read_calc/count[8] ));
   NAND2X1TS \add_x_19_2/U212  (.Y(\add_x_19_2/n166 ), 
	.B(FE_OFN435_offset_6_), 
	.A(\addr_calc/fir_read_calc/count[6] ));
   NAND2X4TS \add_x_19_2/U228  (.Y(\add_x_19_2/n176 ), 
	.B(\addr_calc/fir_read_calc/count[4] ), 
	.A(FE_OFN443_offset_4_));
   NAND2X1TS \add_x_19_2/U237  (.Y(\add_x_19_2/n182 ), 
	.B(FE_OCPN1904_FE_OCPUNCON1066_offset_3_), 
	.A(\addr_calc/fir_read_calc/count[3] ));
   NAND2X1TS \add_x_19_2/U243  (.Y(\add_x_19_2/n185 ), 
	.B(\addr_calc/fir_read_calc/count[2] ), 
	.A(FE_OCPUNCON1065_offset_2_));
   NAND2X1TS \add_x_19_2/U250  (.Y(\add_x_19_2/n189 ), 
	.B(FE_OCP_RBN1974_offset_1_), 
	.A(FE_OFN249_addr_calc_fir_read_calc_count_1_));
   NOR2X2TS \add_x_19_2/U242  (.Y(\add_x_19_2/n184 ), 
	.B(\addr_calc/fir_read_calc/count[2] ), 
	.A(FE_OCPUNCON1065_offset_2_));
   XNOR2X1TS \add_x_19_2/U221  (.Y(\addr_calc/fir_read_addr[4] ), 
	.B(\add_x_19_2/n28 ), 
	.A(\add_x_19_2/n177 ));
   NAND2X1TS \add_x_19_2/U225  (.Y(\add_x_19_2/n28 ), 
	.B(\add_x_19_2/n176 ), 
	.A(\add_x_19_2/n219 ));
   XNOR2X4TS \add_x_19_2/U196  (.Y(\addr_calc/fir_read_addr[7] ), 
	.B(\add_x_19_2/n25 ), 
	.A(\add_x_19_2/n164 ));
   NAND2X1TS \add_x_19_2/U203  (.Y(\add_x_19_2/n25 ), 
	.B(\add_x_19_2/n163 ), 
	.A(\add_x_19_2/n216 ));
   NAND2X1TS \add_x_19_2/U192  (.Y(\add_x_19_2/n24 ), 
	.B(\add_x_19_2/n155 ), 
	.A(\add_x_19_2/n215 ));
   XNOR2X1TS \add_x_19_2/U147  (.Y(\addr_calc/fir_read_addr[13] ), 
	.B(\add_x_19_2/n19 ), 
	.A(\add_x_19_2/n130 ));
   NAND2X1TS \add_x_19_2/U151  (.Y(\add_x_19_2/n19 ), 
	.B(\add_x_19_2/n129 ), 
	.A(\add_x_19_2/n210 ));
   NAND2X2TS \add_x_19_2/U116  (.Y(\add_x_19_2/n15 ), 
	.B(\add_x_19_2/n106 ), 
	.A(\add_x_19_2/n206 ));
   NAND2X1TS \add_x_19_2/U137  (.Y(\add_x_19_2/n17 ), 
	.B(\add_x_19_2/n121 ), 
	.A(\add_x_19_2/n208 ));
   NAND2X1TS \add_x_19_2/U119  (.Y(\add_x_19_2/n106 ), 
	.B(FE_OFN391_offset_17_), 
	.A(\addr_calc/fir_read_calc/count[17] ));
   NAND2X2TS \add_x_19_2/U32  (.Y(\add_x_19_2/n51 ), 
	.B(\add_x_19_2/n53 ), 
	.A(\add_x_19_2/n61 ));
   NAND2X2TS \add_x_19_2/U98  (.Y(\add_x_19_2/n93 ), 
	.B(\add_x_19_2/n95 ), 
	.A(\add_x_19_2/n103 ));
   NAND2X1TS \add_x_19_2/U171  (.Y(\add_x_19_2/n140 ), 
	.B(FE_OCPUNCON652_FE_OFN414_offset_11_), 
	.A(\addr_calc/fir_read_calc/count[11] ));
   NAND2X2TS \add_x_19_2/U133  (.Y(\add_x_19_2/n116 ), 
	.B(\add_x_19_2/n118 ), 
	.A(\add_x_19_2/n126 ));
   NAND2X2TS \add_x_19_2/U164  (.Y(\add_x_19_2/n135 ), 
	.B(\add_x_19_2/n137 ), 
	.A(\add_x_19_2/n149 ));
   NAND2X1TS \add_x_19_2/U220  (.Y(\add_x_19_2/n171 ), 
	.B(FE_OCPUNCON1564_offset_5_), 
	.A(\addr_calc/fir_read_calc/count[5] ));
   NOR2X2TS \add_x_19_1/U236  (.Y(\add_x_19_1/n181 ), 
	.B(FE_OFN447_offset_3_), 
	.A(\addr_calc/fft_write_calc/count[3] ));
   NOR2X4TS \add_x_19_1/U205  (.Y(\add_x_19_1/n162 ), 
	.B(FE_OCP_RBN1842_offset_7_), 
	.A(\addr_calc/fft_write_calc/count[7] ));
   NAND2X6TS \add_x_19_1/U255  (.Y(\add_x_19_1/n191 ), 
	.B(FE_OFN260_addr_calc_fft_write_calc_count_0_), 
	.A(FE_OFN459_offset_0_));
   AOI21X1TS \add_x_19_1/U222  (.Y(\add_x_19_1/n172 ), 
	.B0(\add_x_19_1/n174 ), 
	.A1(\add_x_19_1/n219 ), 
	.A0(\add_x_19_1/n177 ));
   AOI21X4TS \add_x_19_1/U173  (.Y(\add_x_19_1/n141 ), 
	.B0(\add_x_19_1/n143 ), 
	.A1(\add_x_19_1/n213 ), 
	.A0(\add_x_19_1/n146 ));
   OAI21X2TS \add_x_19_1/U181  (.Y(\add_x_19_1/n146 ), 
	.B0(\add_x_19_1/n148 ), 
	.A1(\add_x_19_1/n147 ), 
	.A0(FE_OCP_RBN1956_FE_OFN520_add_x_19_1_n157));
   OAI21X1TS \add_x_19_1/U156  (.Y(\add_x_19_1/n130 ), 
	.B0(\add_x_19_1/n132 ), 
	.A1(\add_x_19_1/n131 ), 
	.A0(\add_x_19_1/n133 ));
   OAI21X1TS \add_x_19_1/U142  (.Y(\add_x_19_1/n122 ), 
	.B0(\add_x_19_1/n124 ), 
	.A1(\add_x_19_1/n123 ), 
	.A0(\add_x_19_1/n125 ));
   AOI21X2TS \add_x_19_1/U148  (.Y(\add_x_19_1/n125 ), 
	.B0(\add_x_19_1/n127 ), 
	.A1(\add_x_19_1/n126 ), 
	.A0(\add_x_19_1/n134 ));
   OAI21X4TS \add_x_19_1/U163  (.Y(\add_x_19_1/n134 ), 
	.B0(\add_x_19_1/n136 ), 
	.A1(\add_x_19_1/n135 ), 
	.A0(FE_OCP_RBN1957_FE_OFN520_add_x_19_1_n157));
   OAI21X2TS \add_x_19_1/U90  (.Y(\add_x_19_1/n88 ), 
	.B0(\add_x_19_1/n90 ), 
	.A1(\add_x_19_1/n89 ), 
	.A0(\add_x_19_1/n91 ));
   OAI21X1TS \add_x_19_1/U31  (.Y(\add_x_19_1/n50 ), 
	.B0(\add_x_19_1/n52 ), 
	.A1(\add_x_19_1/n51 ), 
	.A0(FE_OCP_RBN1379_add_x_19_1_n69));
   OAI21X1TS \add_x_19_1/U55  (.Y(\add_x_19_1/n65 ), 
	.B0(\add_x_19_1/n67 ), 
	.A1(\add_x_19_1/n66 ), 
	.A0(FE_OCP_RBN1379_add_x_19_1_n69));
   NOR2X1TS \add_x_19_1/U10  (.Y(\add_x_19_1/n36 ), 
	.B(FE_OFN341_offset_30_), 
	.A(FE_OFN279_addr_calc_fft_write_calc_count_30_));
   AOI21X2TS \add_x_19_1/U33  (.Y(\add_x_19_1/n52 ), 
	.B0(\add_x_19_1/n54 ), 
	.A1(\add_x_19_1/n62 ), 
	.A0(\add_x_19_1/n53 ));
   OAI21X2TS \add_x_19_1/U35  (.Y(\add_x_19_1/n54 ), 
	.B0(\add_x_19_1/n56 ), 
	.A1(\add_x_19_1/n59 ), 
	.A0(\add_x_19_1/n55 ));
   OAI21X1TS \add_x_19_1/U49  (.Y(\add_x_19_1/n62 ), 
	.B0(\add_x_19_1/n64 ), 
	.A1(\add_x_19_1/n67 ), 
	.A0(\add_x_19_1/n63 ));
   OAI21X2TS \add_x_19_1/U84  (.Y(\add_x_19_1/n85 ), 
	.B0(\add_x_19_1/n87 ), 
	.A1(\add_x_19_1/n90 ), 
	.A0(\add_x_19_1/n86 ));
   OAI21X2TS \add_x_19_1/U101  (.Y(\add_x_19_1/n96 ), 
	.B0(\add_x_19_1/n98 ), 
	.A1(\add_x_19_1/n101 ), 
	.A0(\add_x_19_1/n97 ));
   NOR2X2TS \add_x_19_1/U34  (.Y(\add_x_19_1/n53 ), 
	.B(\add_x_19_1/n55 ), 
	.A(\add_x_19_1/n58 ));
   NOR2X1TS \add_x_19_1/U48  (.Y(\add_x_19_1/n61 ), 
	.B(\add_x_19_1/n63 ), 
	.A(\add_x_19_1/n66 ));
   NOR2X4TS \add_x_19_1/U65  (.Y(\add_x_19_1/n72 ), 
	.B(\add_x_19_1/n74 ), 
	.A(\add_x_19_1/n93 ));
   NOR2X1TS \add_x_19_1/U69  (.Y(\add_x_19_1/n76 ), 
	.B(\add_x_19_1/n78 ), 
	.A(\add_x_19_1/n81 ));
   NOR2X2TS \add_x_19_1/U83  (.Y(\add_x_19_1/n84 ), 
	.B(\add_x_19_1/n86 ), 
	.A(\add_x_19_1/n89 ));
   NOR2X2TS \add_x_19_1/U100  (.Y(\add_x_19_1/n95 ), 
	.B(\add_x_19_1/n97 ), 
	.A(\add_x_19_1/n100 ));
   OAI21X1TS \add_x_19_1/U150  (.Y(\add_x_19_1/n127 ), 
	.B0(\add_x_19_1/n129 ), 
	.A1(\add_x_19_1/n132 ), 
	.A0(\add_x_19_1/n128 ));
   NOR2X1TS \add_x_19_1/U139  (.Y(\add_x_19_1/n120 ), 
	.B(\addr_calc/fft_write_calc/count[15] ), 
	.A(FE_OFN399_offset_15_));
   NOR2X2TS \add_x_19_1/U149  (.Y(\add_x_19_1/n126 ), 
	.B(\add_x_19_1/n131 ), 
	.A(\add_x_19_1/n128 ));
   NOR2X2TS \add_x_19_1/U184  (.Y(\add_x_19_1/n149 ), 
	.B(\add_x_19_1/n151 ), 
	.A(\add_x_19_1/n154 ));
   NOR2X1TS \add_x_19_1/U249  (.Y(\add_x_19_1/n188 ), 
	.B(\addr_calc/fft_write_calc/count[1] ), 
	.A(FE_OCP_RBN1973_offset_1_));
   XOR2X1TS \add_x_19_1/U213  (.Y(\addr_calc/fft_write_addr[5] ), 
	.B(\add_x_19_1/n27 ), 
	.A(\add_x_19_1/n172 ));
   XOR2X4TS \add_x_19_1/U161  (.Y(\addr_calc/fft_write_addr[11] ), 
	.B(\add_x_19_1/n21 ), 
	.A(\add_x_19_1/n141 ));
   NAND2X1TS \add_x_19_1/U11  (.Y(\add_x_19_1/n37 ), 
	.B(FE_OFN341_offset_30_), 
	.A(FE_OFN279_addr_calc_fft_write_calc_count_30_));
   NAND2X1TS \add_x_19_1/U19  (.Y(\add_x_19_1/n42 ), 
	.B(FE_OFN345_offset_29_), 
	.A(\addr_calc/fft_write_calc/count[29] ));
   NAND2X1TS \add_x_19_1/U29  (.Y(\add_x_19_1/n49 ), 
	.B(FE_OFN349_offset_28_), 
	.A(n2557));
   NAND2X1TS \add_x_19_1/U39  (.Y(\add_x_19_1/n56 ), 
	.B(FE_OFN353_offset_27_), 
	.A(n1913));
   NAND2X1TS \add_x_19_1/U45  (.Y(\add_x_19_1/n59 ), 
	.B(FE_OFN358_offset_26_), 
	.A(\addr_calc/fft_write_calc/count[26] ));
   NAND2X1TS \add_x_19_1/U53  (.Y(\add_x_19_1/n64 ), 
	.B(FE_OFN361_offset_25_), 
	.A(n1915));
   NAND2X1TS \add_x_19_1/U74  (.Y(\add_x_19_1/n79 ), 
	.B(FE_OCPUNCON1069_FE_OFN369_offset_23_), 
	.A(\addr_calc/fft_write_calc/count[23] ));
   NAND2X1TS \add_x_19_1/U80  (.Y(\add_x_19_1/n82 ), 
	.B(FE_OFN374_offset_22_), 
	.A(FE_OFN284_addr_calc_fft_write_calc_count_22_));
   NAND2X1TS \add_x_19_1/U88  (.Y(\add_x_19_1/n87 ), 
	.B(FE_OFN377_offset_21_), 
	.A(n1918));
   NAND2X1TS \add_x_19_1/U94  (.Y(\add_x_19_1/n90 ), 
	.B(FE_OFN557_n2441), 
	.A(FE_OFN281_addr_calc_fft_write_calc_count_20_));
   NAND2X1TS \add_x_19_1/U105  (.Y(\add_x_19_1/n98 ), 
	.B(FE_OFN382_offset_19_), 
	.A(n1922));
   NAND2X1TS \add_x_19_1/U111  (.Y(\add_x_19_1/n101 ), 
	.B(FE_OFN386_offset_18_), 
	.A(n2020));
   NAND2X1TS \add_x_19_1/U119  (.Y(\add_x_19_1/n106 ), 
	.B(FE_OFN390_offset_17_), 
	.A(\addr_calc/fft_write_calc/count[17] ));
   NOR2X1TS \add_x_19_1/U52  (.Y(\add_x_19_1/n63 ), 
	.B(FE_OFN361_offset_25_), 
	.A(n1915));
   NOR2X1TS \add_x_19_1/U58  (.Y(\add_x_19_1/n66 ), 
	.B(FE_OFN365_offset_24_), 
	.A(FE_OFN277_addr_calc_fft_write_calc_count_24_));
   NOR2X1TS \add_x_19_1/U79  (.Y(\add_x_19_1/n81 ), 
	.B(FE_OFN374_offset_22_), 
	.A(FE_OFN284_addr_calc_fft_write_calc_count_22_));
   NOR2X1TS \add_x_19_1/U87  (.Y(\add_x_19_1/n86 ), 
	.B(FE_OFN377_offset_21_), 
	.A(n1918));
   NOR2X1TS \add_x_19_1/U93  (.Y(\add_x_19_1/n89 ), 
	.B(FE_OFN557_n2441), 
	.A(FE_OFN281_addr_calc_fft_write_calc_count_20_));
   NOR2X1TS \add_x_19_1/U104  (.Y(\add_x_19_1/n97 ), 
	.B(FE_OFN382_offset_19_), 
	.A(n1922));
   NOR2X1TS \add_x_19_1/U110  (.Y(\add_x_19_1/n100 ), 
	.B(FE_OFN386_offset_18_), 
	.A(n2020));
   NOR2X1TS \add_x_19_1/U118  (.Y(\add_x_19_1/n105 ), 
	.B(FE_OFN390_offset_17_), 
	.A(\addr_calc/fft_write_calc/count[17] ));
   NAND2X1TS \add_x_19_1/U140  (.Y(\add_x_19_1/n121 ), 
	.B(FE_OFN399_offset_15_), 
	.A(\addr_calc/fft_write_calc/count[15] ));
   NAND2X1TS \add_x_19_1/U146  (.Y(\add_x_19_1/n124 ), 
	.B(FE_OFN403_offset_14_), 
	.A(FE_OFN259_addr_calc_fft_write_calc_count_14_));
   NAND2X1TS \add_x_19_1/U154  (.Y(\add_x_19_1/n129 ), 
	.B(FE_OCPUNCON1941_offset_13_), 
	.A(\addr_calc/fft_write_calc/count[13] ));
   NAND2X1TS \add_x_19_1/U160  (.Y(\add_x_19_1/n132 ), 
	.B(FE_OFN410_offset_12_), 
	.A(\addr_calc/fft_write_calc/count[12] ));
   NAND2X1TS \add_x_19_1/U179  (.Y(\add_x_19_1/n145 ), 
	.B(FE_OFN418_offset_10_), 
	.A(\addr_calc/fft_write_calc/count[10] ));
   NAND2X1TS \add_x_19_1/U189  (.Y(\add_x_19_1/n152 ), 
	.B(FE_OFN422_offset_9_), 
	.A(\addr_calc/fft_write_calc/count[9] ));
   NOR2X1TS \add_x_19_1/U153  (.Y(\add_x_19_1/n128 ), 
	.B(FE_OCPUNCON1941_offset_13_), 
	.A(\addr_calc/fft_write_calc/count[13] ));
   NOR2X1TS \add_x_19_1/U159  (.Y(\add_x_19_1/n131 ), 
	.B(FE_OFN410_offset_12_), 
	.A(\addr_calc/fft_write_calc/count[12] ));
   NOR2X1TS \add_x_19_1/U194  (.Y(\add_x_19_1/n154 ), 
	.B(FE_OFN427_offset_8_), 
	.A(\addr_calc/fft_write_calc/count[8] ));
   NAND2X1TS \add_x_19_1/U206  (.Y(\add_x_19_1/n163 ), 
	.B(FE_OCP_RBN1842_offset_7_), 
	.A(\addr_calc/fft_write_calc/count[7] ));
   NAND2X1TS \add_x_19_1/U212  (.Y(\add_x_19_1/n166 ), 
	.B(FE_OCPUNCON1684_offset_6_), 
	.A(FE_OFN271_addr_calc_fft_write_calc_count_6_));
   NOR2X2TS \add_x_19_1/U227  (.Y(\add_x_19_1/n175 ), 
	.B(\addr_calc/fft_write_calc/count[4] ), 
	.A(FE_OCPUNCON1875_offset_4_));
   NAND2X1TS \add_x_19_1/U237  (.Y(\add_x_19_1/n182 ), 
	.B(FE_OFN447_offset_3_), 
	.A(\addr_calc/fft_write_calc/count[3] ));
   NAND2X6TS \add_x_19_1/U243  (.Y(\add_x_19_1/n185 ), 
	.B(\addr_calc/fft_write_calc/count[2] ), 
	.A(FE_OFN451_offset_2_));
   NAND2X1TS \add_x_19_1/U250  (.Y(\add_x_19_1/n189 ), 
	.B(\addr_calc/fft_write_calc/count[1] ), 
	.A(FE_OCP_RBN1973_offset_1_));
   NOR2X1TS \add_x_19_1/U242  (.Y(\add_x_19_1/n184 ), 
	.B(\addr_calc/fft_write_calc/count[2] ), 
	.A(FE_OFN451_offset_2_));
   XNOR2X1TS \add_x_19_1/U221  (.Y(\addr_calc/fft_write_addr[4] ), 
	.B(\add_x_19_1/n28 ), 
	.A(\add_x_19_1/n177 ));
   NAND2X1TS \add_x_19_1/U225  (.Y(\add_x_19_1/n28 ), 
	.B(\add_x_19_1/n176 ), 
	.A(\add_x_19_1/n219 ));
   NAND2X2TS \add_x_19_1/U168  (.Y(\add_x_19_1/n21 ), 
	.B(\add_x_19_1/n140 ), 
	.A(\add_x_19_1/n212 ));
   XNOR2X2TS \add_x_19_1/U147  (.Y(\addr_calc/fft_write_addr[13] ), 
	.B(\add_x_19_1/n19 ), 
	.A(\add_x_19_1/n130 ));
   NAND2X1TS \add_x_19_1/U151  (.Y(\add_x_19_1/n19 ), 
	.B(\add_x_19_1/n129 ), 
	.A(\add_x_19_1/n210 ));
   NAND2X1TS \add_x_19_1/U137  (.Y(\add_x_19_1/n17 ), 
	.B(\add_x_19_1/n121 ), 
	.A(\add_x_19_1/n208 ));
   XNOR2X4TS \add_x_19_1/U12  (.Y(\addr_calc/fft_write_addr[29] ), 
	.B(\add_x_19_1/n43 ), 
	.A(\add_x_19_1/n3 ));
   NAND2X1TS \add_x_19_1/U16  (.Y(\add_x_19_1/n3 ), 
	.B(\add_x_19_1/n42 ), 
	.A(n2632));
   NAND2X2TS \add_x_19_1/U85  (.Y(\add_x_19_1/n11 ), 
	.B(\add_x_19_1/n87 ), 
	.A(\add_x_19_1/n202 ));
   NAND2X1TS \add_x_19_1/U26  (.Y(\add_x_19_1/n4 ), 
	.B(\add_x_19_1/n49 ), 
	.A(\add_x_19_1/n195 ));
   NAND2X1TS \add_x_19_1/U50  (.Y(\add_x_19_1/n7 ), 
	.B(\add_x_19_1/n64 ), 
	.A(\add_x_19_1/n198 ));
   NAND2X1TS \add_x_19_1/U32  (.Y(\add_x_19_1/n51 ), 
	.B(\add_x_19_1/n53 ), 
	.A(\add_x_19_1/n61 ));
   NAND2X2TS \add_x_19_1/U67  (.Y(\add_x_19_1/n74 ), 
	.B(\add_x_19_1/n76 ), 
	.A(\add_x_19_1/n84 ));
   NAND2X4TS \add_x_19_1/U98  (.Y(\add_x_19_1/n93 ), 
	.B(\add_x_19_1/n95 ), 
	.A(\add_x_19_1/n103 ));
   NAND2X1TS \add_x_19_1/U171  (.Y(\add_x_19_1/n140 ), 
	.B(FE_OCPN1905_FE_OCPUNCON1873_offset_11_), 
	.A(n1667));
   NAND2X1TS \add_x_19_1/U133  (.Y(\add_x_19_1/n116 ), 
	.B(\add_x_19_1/n126 ), 
	.A(\add_x_19_1/n118 ));
   NAND2X4TS \add_x_19_1/U164  (.Y(\add_x_19_1/n135 ), 
	.B(\add_x_19_1/n137 ), 
	.A(\add_x_19_1/n149 ));
   NOR2X2TS \add_x_19_3/U118  (.Y(\add_x_19_3/n105 ), 
	.B(FE_OFN393_offset_17_), 
	.A(n1886));
   NOR2X8TS \add_x_19_3/U219  (.Y(\add_x_19_3/n170 ), 
	.B(FE_OCP_RBN1495_offset_5_), 
	.A(\addr_calc/fir_write_calc/count[5] ));
   OAI21X2TS \add_x_19_3/U70  (.Y(\add_x_19_3/n77 ), 
	.B0(\add_x_19_3/n79 ), 
	.A1(\add_x_19_3/n82 ), 
	.A0(\add_x_19_3/n78 ));
   XOR2X2TS \add_x_19_3/U238  (.Y(\addr_calc/fir_write_addr[2] ), 
	.B(\add_x_19_3/n30 ), 
	.A(\add_x_19_3/n186 ));
   AOI21X1TS \add_x_19_3/U222  (.Y(\add_x_19_3/n172 ), 
	.B0(\add_x_19_3/n174 ), 
	.A1(\add_x_19_3/n219 ), 
	.A0(\add_x_19_3/n177 ));
   AOI21X2TS \add_x_19_3/U214  (.Y(\add_x_19_3/n167 ), 
	.B0(\add_x_19_3/n169 ), 
	.A1(\add_x_19_3/n168 ), 
	.A0(\add_x_19_3/n177 ));
   XOR2X1TS \add_x_19_3/U190  (.Y(\addr_calc/fir_write_addr[8] ), 
	.B(\add_x_19_3/n24 ), 
	.A(\add_x_19_3/n156 ));
   OAI21X1TS \add_x_19_3/U142  (.Y(\add_x_19_3/n122 ), 
	.B0(\add_x_19_3/n124 ), 
	.A1(\add_x_19_3/n123 ), 
	.A0(\add_x_19_3/n125 ));
   AOI21X4TS \add_x_19_3/U148  (.Y(\add_x_19_3/n125 ), 
	.B0(\add_x_19_3/n127 ), 
	.A1(\add_x_19_3/n126 ), 
	.A0(\add_x_19_3/n134 ));
   OAI21X1TS \add_x_19_3/U107  (.Y(\add_x_19_3/n99 ), 
	.B0(\add_x_19_3/n101 ), 
	.A1(\add_x_19_3/n100 ), 
	.A0(\add_x_19_3/n102 ));
   AOI21X4TS \add_x_19_3/U113  (.Y(\add_x_19_3/n102 ), 
	.B0(\add_x_19_3/n104 ), 
	.A1(\add_x_19_3/n103 ), 
	.A0(FE_OCP_RBN1378_add_x_19_3_n113));
   OAI21X2TS \add_x_19_3/U90  (.Y(\add_x_19_3/n88 ), 
	.B0(\add_x_19_3/n90 ), 
	.A1(\add_x_19_3/n89 ), 
	.A0(FE_OCP_RBN1381_add_x_19_3_n92));
   NOR2X1TS \add_x_19_3/U10  (.Y(\add_x_19_3/n36 ), 
	.B(FE_OFN344_offset_30_), 
	.A(\addr_calc/fir_write_calc/count[30] ));
   OAI21X2TS \add_x_19_3/U25  (.Y(\add_x_19_3/n47 ), 
	.B0(\add_x_19_3/n49 ), 
	.A1(\add_x_19_3/n48 ), 
	.A0(\add_x_19_3/n52 ));
   OAI21X1TS \add_x_19_3/U35  (.Y(\add_x_19_3/n54 ), 
	.B0(\add_x_19_3/n56 ), 
	.A1(\add_x_19_3/n59 ), 
	.A0(\add_x_19_3/n55 ));
   NOR2X2TS \add_x_19_3/U28  (.Y(\add_x_19_3/n48 ), 
	.B(FE_OFN352_offset_28_), 
	.A(\addr_calc/fir_write_calc/count[28] ));
   OAI21X2TS \add_x_19_3/U49  (.Y(\add_x_19_3/n62 ), 
	.B0(\add_x_19_3/n64 ), 
	.A1(\add_x_19_3/n67 ), 
	.A0(\add_x_19_3/n63 ));
   NOR2X2TS \add_x_19_3/U48  (.Y(\add_x_19_3/n61 ), 
	.B(\add_x_19_3/n63 ), 
	.A(\add_x_19_3/n66 ));
   AOI21X2TS \add_x_19_3/U68  (.Y(\add_x_19_3/n75 ), 
	.B0(\add_x_19_3/n77 ), 
	.A1(\add_x_19_3/n85 ), 
	.A0(\add_x_19_3/n76 ));
   OAI21X1TS \add_x_19_3/U84  (.Y(\add_x_19_3/n85 ), 
	.B0(\add_x_19_3/n87 ), 
	.A1(\add_x_19_3/n90 ), 
	.A0(\add_x_19_3/n86 ));
   NOR2X4TS \add_x_19_3/U69  (.Y(\add_x_19_3/n76 ), 
	.B(\add_x_19_3/n78 ), 
	.A(\add_x_19_3/n81 ));
   NOR2X4TS \add_x_19_3/U83  (.Y(\add_x_19_3/n84 ), 
	.B(\add_x_19_3/n86 ), 
	.A(\add_x_19_3/n89 ));
   NOR2X4TS \add_x_19_3/U100  (.Y(\add_x_19_3/n95 ), 
	.B(\add_x_19_3/n97 ), 
	.A(\add_x_19_3/n100 ));
   NOR2X4TS \add_x_19_3/U114  (.Y(\add_x_19_3/n103 ), 
	.B(\add_x_19_3/n105 ), 
	.A(\add_x_19_3/n110 ));
   NOR2X4TS \add_x_19_3/U166  (.Y(\add_x_19_3/n137 ), 
	.B(\add_x_19_3/n144 ), 
	.A(\add_x_19_3/n139 ));
   NOR2X8TS \add_x_19_3/U170  (.Y(\add_x_19_3/n139 ), 
	.B(\addr_calc/fir_write_calc/count[11] ), 
	.A(FE_OCPUNCON656_FE_OFN414_offset_11_));
   NOR2X1TS \add_x_19_3/U184  (.Y(\add_x_19_3/n149 ), 
	.B(\add_x_19_3/n154 ), 
	.A(\add_x_19_3/n151 ));
   NOR2X6TS \add_x_19_3/U215  (.Y(\add_x_19_3/n168 ), 
	.B(\add_x_19_3/n170 ), 
	.A(\add_x_19_3/n175 ));
   NOR2X2TS \add_x_19_3/U249  (.Y(\add_x_19_3/n188 ), 
	.B(FE_OCPUNCON1874_offset_1_), 
	.A(FE_OFN242_addr_calc_fir_write_calc_count_1_));
   XOR2X2TS \add_x_19_3/U213  (.Y(\addr_calc/fir_write_addr[5] ), 
	.B(\add_x_19_3/n27 ), 
	.A(\add_x_19_3/n172 ));
   CLKXOR2X2TS \add_x_19_3/U207  (.Y(\addr_calc/fir_write_addr[6] ), 
	.B(\add_x_19_3/n26 ), 
	.A(\add_x_19_3/n167 ));
   XOR2X4TS \add_x_19_3/U141  (.Y(\addr_calc/fir_write_addr[14] ), 
	.B(\add_x_19_3/n18 ), 
	.A(\add_x_19_3/n125 ));
   NAND2X1TS \add_x_19_3/U11  (.Y(\add_x_19_3/n37 ), 
	.B(FE_OFN344_offset_30_), 
	.A(\addr_calc/fir_write_calc/count[30] ));
   NAND2X1TS \add_x_19_3/U19  (.Y(\add_x_19_3/n42 ), 
	.B(FE_OFN348_offset_29_), 
	.A(FE_OFN273_addr_calc_fir_write_calc_count_29_));
   NAND2X1TS \add_x_19_3/U29  (.Y(\add_x_19_3/n49 ), 
	.B(FE_OFN352_offset_28_), 
	.A(n1896));
   NAND2X1TS \add_x_19_3/U39  (.Y(\add_x_19_3/n56 ), 
	.B(FE_OFN356_offset_27_), 
	.A(n1835));
   NAND2X1TS \add_x_19_3/U45  (.Y(\add_x_19_3/n59 ), 
	.B(FE_OFN359_offset_26_), 
	.A(FE_OFN267_addr_calc_fir_write_calc_count_26_));
   NAND2X1TS \add_x_19_3/U53  (.Y(\add_x_19_3/n64 ), 
	.B(FE_OFN363_offset_25_), 
	.A(FE_OFN231_addr_calc_fir_write_calc_count_25_));
   NAND2X2TS \add_x_19_3/U59  (.Y(\add_x_19_3/n67 ), 
	.B(FE_OFN368_offset_24_), 
	.A(\addr_calc/fir_write_calc/count[24] ));
   NAND2X1TS \add_x_19_3/U74  (.Y(\add_x_19_3/n79 ), 
	.B(FE_OFN371_offset_23_), 
	.A(\addr_calc/fir_write_calc/count[23] ));
   NAND2X1TS \add_x_19_3/U80  (.Y(\add_x_19_3/n82 ), 
	.B(FE_OFN375_offset_22_), 
	.A(\addr_calc/fir_write_calc/count[22] ));
   NAND2X1TS \add_x_19_3/U88  (.Y(\add_x_19_3/n87 ), 
	.B(FE_OCPUNCON1078_FE_OFN377_offset_21_), 
	.A(n1892));
   NAND2X2TS \add_x_19_3/U94  (.Y(\add_x_19_3/n90 ), 
	.B(n2441), 
	.A(FE_OFN283_addr_calc_fir_write_calc_count_20_));
   NAND2X1TS \add_x_19_3/U105  (.Y(\add_x_19_3/n98 ), 
	.B(FE_OCPUNCON1079_FE_OFN382_offset_19_), 
	.A(n1670));
   NAND2X1TS \add_x_19_3/U111  (.Y(\add_x_19_3/n101 ), 
	.B(FE_OCPUNCON1080_FE_OFN386_offset_18_), 
	.A(\addr_calc/fir_write_calc/count[18] ));
   NOR2X4TS \add_x_19_3/U79  (.Y(\add_x_19_3/n81 ), 
	.B(FE_OFN375_offset_22_), 
	.A(n1668));
   NOR2X1TS \add_x_19_3/U93  (.Y(\add_x_19_3/n89 ), 
	.B(n2441), 
	.A(FE_OFN283_addr_calc_fir_write_calc_count_20_));
   NOR2X1TS \add_x_19_3/U110  (.Y(\add_x_19_3/n100 ), 
	.B(n2006), 
	.A(FE_OCPUNCON1080_FE_OFN386_offset_18_));
   NAND2X2TS \add_x_19_3/U140  (.Y(\add_x_19_3/n121 ), 
	.B(FE_OFN400_offset_15_), 
	.A(n1883));
   NAND2X2TS \add_x_19_3/U146  (.Y(\add_x_19_3/n124 ), 
	.B(FE_OFN404_offset_14_), 
	.A(n2003));
   NAND2X2TS \add_x_19_3/U154  (.Y(\add_x_19_3/n129 ), 
	.B(FE_OCPUNCON1943_FE_OFN407_offset_13_), 
	.A(\addr_calc/fir_write_calc/count[13] ));
   NAND2X4TS \add_x_19_3/U179  (.Y(\add_x_19_3/n145 ), 
	.B(FE_OCPUNCON657_FE_OFN418_offset_10_), 
	.A(\addr_calc/fir_write_calc/count[10] ));
   NAND2X2TS \add_x_19_3/U189  (.Y(\add_x_19_3/n152 ), 
	.B(FE_OCPUNCON658_FE_OFN422_offset_9_), 
	.A(\addr_calc/fir_write_calc/count[9] ));
   NOR2X8TS \add_x_19_3/U153  (.Y(\add_x_19_3/n128 ), 
	.B(FE_OCPUNCON1943_FE_OFN407_offset_13_), 
	.A(\addr_calc/fir_write_calc/count[13] ));
   NOR2X6TS \add_x_19_3/U178  (.Y(\add_x_19_3/n144 ), 
	.B(FE_OCPUNCON657_FE_OFN418_offset_10_), 
	.A(\addr_calc/fir_write_calc/count[10] ));
   NOR2X4TS \add_x_19_3/U188  (.Y(\add_x_19_3/n151 ), 
	.B(\addr_calc/fir_write_calc/count[9] ), 
	.A(FE_OCPUNCON658_FE_OFN422_offset_9_));
   NOR2X4TS \add_x_19_3/U194  (.Y(\add_x_19_3/n154 ), 
	.B(FE_OFN428_offset_8_), 
	.A(FE_OFN255_addr_calc_fir_write_calc_count_8_));
   NAND2X6TS \add_x_19_3/U206  (.Y(\add_x_19_3/n163 ), 
	.B(\addr_calc/fir_write_calc/count[7] ), 
	.A(FE_OCPUNCON1278_offset_7_));
   NAND2X1TS \add_x_19_3/U212  (.Y(\add_x_19_3/n166 ), 
	.B(FE_OCPUNCON726_FE_OFN435_offset_6_), 
	.A(FE_OFN253_addr_calc_fir_write_calc_count_6_));
   NAND2X2TS \add_x_19_3/U228  (.Y(\add_x_19_3/n176 ), 
	.B(FE_OFN241_addr_calc_fir_write_calc_count_4_), 
	.A(FE_OCPUNCON1425_FE_OFN443_offset_4_));
   NOR2X6TS \add_x_19_3/U227  (.Y(\add_x_19_3/n175 ), 
	.B(FE_OFN241_addr_calc_fir_write_calc_count_4_), 
	.A(FE_OCPN1224_FE_OFN445_offset_4_));
   NAND2X4TS \add_x_19_3/U237  (.Y(\add_x_19_3/n182 ), 
	.B(FE_OFN449_offset_3_), 
	.A(\addr_calc/fir_write_calc/count[3] ));
   NAND2X1TS \add_x_19_3/U250  (.Y(\add_x_19_3/n189 ), 
	.B(FE_OFN242_addr_calc_fir_write_calc_count_1_), 
	.A(FE_OCPUNCON1874_offset_1_));
   NAND2X1TS \add_x_19_3/U240  (.Y(\add_x_19_3/n30 ), 
	.B(\add_x_19_3/n185 ), 
	.A(\add_x_19_3/n221 ));
   XNOR2XLTS \add_x_19_3/U221  (.Y(\addr_calc/fir_write_addr[4] ), 
	.B(\add_x_19_3/n28 ), 
	.A(\add_x_19_3/n177 ));
   NAND2X1TS \add_x_19_3/U225  (.Y(\add_x_19_3/n28 ), 
	.B(\add_x_19_3/n176 ), 
	.A(\add_x_19_3/n219 ));
   NAND2X1TS \add_x_19_3/U217  (.Y(\add_x_19_3/n27 ), 
	.B(\add_x_19_3/n171 ), 
	.A(\add_x_19_3/n218 ));
   NAND2X1TS \add_x_19_3/U209  (.Y(\add_x_19_3/n26 ), 
	.B(\add_x_19_3/n166 ), 
	.A(\add_x_19_3/n217 ));
   NAND2X1TS \add_x_19_3/U192  (.Y(\add_x_19_3/n24 ), 
	.B(\add_x_19_3/n155 ), 
	.A(\add_x_19_3/n215 ));
   XNOR2X2TS \add_x_19_3/U172  (.Y(\addr_calc/fir_write_addr[10] ), 
	.B(\add_x_19_3/n22 ), 
	.A(\add_x_19_3/n146 ));
   NAND2X1TS \add_x_19_3/U176  (.Y(\add_x_19_3/n22 ), 
	.B(\add_x_19_3/n145 ), 
	.A(\add_x_19_3/n213 ));
   NAND2XLTS \add_x_19_3/U143  (.Y(\add_x_19_3/n18 ), 
	.B(\add_x_19_3/n124 ), 
	.A(n1545));
   XNOR2X4TS \add_x_19_3/U128  (.Y(\addr_calc/fir_write_addr[15] ), 
	.B(\add_x_19_3/n17 ), 
	.A(\add_x_19_3/n122 ));
   NAND2X1TS \add_x_19_3/U137  (.Y(\add_x_19_3/n17 ), 
	.B(\add_x_19_3/n121 ), 
	.A(\add_x_19_3/n208 ));
   XNOR2X4TS \add_x_19_3/U95  (.Y(\addr_calc/fir_write_addr[19] ), 
	.B(\add_x_19_3/n13 ), 
	.A(\add_x_19_3/n99 ));
   NAND2X1TS \add_x_19_3/U102  (.Y(\add_x_19_3/n13 ), 
	.B(\add_x_19_3/n98 ), 
	.A(\add_x_19_3/n204 ));
   XNOR2X2TS \add_x_19_3/U81  (.Y(\addr_calc/fir_write_addr[21] ), 
	.B(\add_x_19_3/n11 ), 
	.A(\add_x_19_3/n88 ));
   NAND2X2TS \add_x_19_3/U85  (.Y(\add_x_19_3/n11 ), 
	.B(\add_x_19_3/n87 ), 
	.A(\add_x_19_3/n202 ));
   NAND2X1TS \add_x_19_3/U26  (.Y(\add_x_19_3/n4 ), 
	.B(\add_x_19_3/n49 ), 
	.A(\add_x_19_3/n195 ));
   XNOR2X4TS \add_x_19_3/U46  (.Y(\addr_calc/fir_write_addr[25] ), 
	.B(\add_x_19_3/n7 ), 
	.A(\add_x_19_3/n65 ));
   NAND2X2TS \add_x_19_3/U50  (.Y(\add_x_19_3/n7 ), 
	.B(\add_x_19_3/n64 ), 
	.A(\add_x_19_3/n198 ));
   NAND2X1TS \add_x_19_3/U119  (.Y(\add_x_19_3/n106 ), 
	.B(FE_OFN393_offset_17_), 
	.A(n1886));
   NAND2X2TS \add_x_19_3/U67  (.Y(\add_x_19_3/n74 ), 
	.B(\add_x_19_3/n76 ), 
	.A(\add_x_19_3/n84 ));
   NAND2X2TS \add_x_19_3/U171  (.Y(\add_x_19_3/n140 ), 
	.B(\addr_calc/fir_write_calc/count[11] ), 
	.A(FE_OCPUNCON656_FE_OFN414_offset_11_));
   NAND2X2TS \add_x_19_3/U164  (.Y(\add_x_19_3/n135 ), 
	.B(\add_x_19_3/n137 ), 
	.A(\add_x_19_3/n149 ));
   NAND2X1TS \add_x_19_3/U220  (.Y(\add_x_19_3/n171 ), 
	.B(FE_OCP_RBN1495_offset_5_), 
	.A(\addr_calc/fir_write_calc/count[5] ));
   NOR2X4TS \add_x_19_5/U236  (.Y(\add_x_19_5/n181 ), 
	.B(FE_OFN250_addr_calc_iir_write_calc_count_3_), 
	.A(FE_OCPUNCON1075_FE_OFN447_offset_3_));
   NAND2X4TS \add_x_19_5/U255  (.Y(\add_x_19_5/n191 ), 
	.B(FE_OCPUNCON1077_FE_OFN459_offset_0_), 
	.A(\addr_calc/iir_write_calc/count[0] ));
   XOR2X1TS \add_x_19_5/U244  (.Y(\addr_calc/iir_write_addr[1] ), 
	.B(\add_x_19_5/n191 ), 
	.A(\add_x_19_5/n31 ));
   AOI21X2TS \add_x_19_5/U214  (.Y(\add_x_19_5/n167 ), 
	.B0(\add_x_19_5/n169 ), 
	.A1(\add_x_19_5/n168 ), 
	.A0(n1818));
   OAI21X1TS \add_x_19_5/U191  (.Y(\add_x_19_5/n153 ), 
	.B0(\add_x_19_5/n155 ), 
	.A1(\add_x_19_5/n154 ), 
	.A0(\add_x_19_5/n156 ));
   OAI21X4TS \add_x_19_5/U181  (.Y(\add_x_19_5/n146 ), 
	.B0(\add_x_19_5/n148 ), 
	.A1(\add_x_19_5/n147 ), 
	.A0(\add_x_19_5/n156 ));
   AOI21X2TS \add_x_19_5/U121  (.Y(\add_x_19_5/n107 ), 
	.B0(\add_x_19_5/n109 ), 
	.A1(\add_x_19_5/n207 ), 
	.A0(\add_x_19_5/n112 ));
   OAI21X4TS \add_x_19_5/U31  (.Y(\add_x_19_5/n50 ), 
	.B0(\add_x_19_5/n52 ), 
	.A1(\add_x_19_5/n51 ), 
	.A0(\add_x_19_5/n68 ));
   OAI21X1TS \add_x_19_5/U55  (.Y(\add_x_19_5/n65 ), 
	.B0(\add_x_19_5/n67 ), 
	.A1(\add_x_19_5/n66 ), 
	.A0(\add_x_19_5/n68 ));
   NOR2X1TS \add_x_19_5/U10  (.Y(\add_x_19_5/n36 ), 
	.B(FE_OFN559_offset_30_), 
	.A(FE_OFN239_addr_calc_iir_write_calc_count_30_));
   OAI21X2TS \add_x_19_5/U49  (.Y(\add_x_19_5/n62 ), 
	.B0(\add_x_19_5/n64 ), 
	.A1(\add_x_19_5/n67 ), 
	.A0(\add_x_19_5/n63 ));
   OAI21X2TS \add_x_19_5/U101  (.Y(\add_x_19_5/n96 ), 
	.B0(\add_x_19_5/n98 ), 
	.A1(\add_x_19_5/n101 ), 
	.A0(\add_x_19_5/n97 ));
   NOR2X2TS \add_x_19_5/U28  (.Y(\add_x_19_5/n48 ), 
	.B(FE_OFN351_offset_28_), 
	.A(n1974));
   NOR2X2TS \add_x_19_5/U34  (.Y(\add_x_19_5/n53 ), 
	.B(\add_x_19_5/n55 ), 
	.A(\add_x_19_5/n58 ));
   NOR2X2TS \add_x_19_5/U48  (.Y(\add_x_19_5/n61 ), 
	.B(\add_x_19_5/n63 ), 
	.A(\add_x_19_5/n66 ));
   NOR2X4TS \add_x_19_5/U65  (.Y(\add_x_19_5/n72 ), 
	.B(\add_x_19_5/n74 ), 
	.A(\add_x_19_5/n93 ));
   NOR2X2TS \add_x_19_5/U83  (.Y(\add_x_19_5/n84 ), 
	.B(\add_x_19_5/n86 ), 
	.A(\add_x_19_5/n89 ));
   NOR2X2TS \add_x_19_5/U100  (.Y(\add_x_19_5/n95 ), 
	.B(\add_x_19_5/n97 ), 
	.A(\add_x_19_5/n100 ));
   OAI21X4TS \add_x_19_5/U150  (.Y(\add_x_19_5/n127 ), 
	.B0(\add_x_19_5/n129 ), 
	.A1(\add_x_19_5/n132 ), 
	.A0(\add_x_19_5/n128 ));
   NOR2X4TS \add_x_19_5/U139  (.Y(\add_x_19_5/n120 ), 
	.B(FE_OFN229_addr_calc_iir_write_calc_count_15_), 
	.A(FE_OCPUNCON1942_FE_OFN399_offset_15_));
   NOR2X2TS \add_x_19_5/U149  (.Y(\add_x_19_5/n126 ), 
	.B(\add_x_19_5/n128 ), 
	.A(\add_x_19_5/n131 ));
   NOR2X2TS \add_x_19_5/U166  (.Y(\add_x_19_5/n137 ), 
	.B(\add_x_19_5/n144 ), 
	.A(\add_x_19_5/n139 ));
   NOR2X8TS \add_x_19_5/U170  (.Y(\add_x_19_5/n139 ), 
	.B(FE_OFN417_offset_11_), 
	.A(\addr_calc/iir_write_calc/count[11] ));
   NOR2X2TS \add_x_19_5/U184  (.Y(\add_x_19_5/n149 ), 
	.B(\add_x_19_5/n151 ), 
	.A(\add_x_19_5/n154 ));
   OAI21X4TS \add_x_19_5/U216  (.Y(\add_x_19_5/n169 ), 
	.B0(\add_x_19_5/n171 ), 
	.A1(\add_x_19_5/n176 ), 
	.A0(\add_x_19_5/n170 ));
   NOR2X4TS \add_x_19_5/U201  (.Y(\add_x_19_5/n160 ), 
	.B(\add_x_19_5/n165 ), 
	.A(\add_x_19_5/n162 ));
   NOR2X2TS \add_x_19_5/U215  (.Y(\add_x_19_5/n168 ), 
	.B(\add_x_19_5/n175 ), 
	.A(\add_x_19_5/n170 ));
   OAI21X4TS \add_x_19_5/U246  (.Y(\add_x_19_5/n187 ), 
	.B0(\add_x_19_5/n189 ), 
	.A1(\add_x_19_5/n188 ), 
	.A0(\add_x_19_5/n191 ));
   NOR2X8TS \add_x_19_5/U249  (.Y(\add_x_19_5/n188 ), 
	.B(\addr_calc/iir_write_calc/count[1] ), 
	.A(FE_OCP_RBN1919_offset_1_));
   NOR2X2TS \add_x_19_5/U232  (.Y(\add_x_19_5/n179 ), 
	.B(\add_x_19_5/n181 ), 
	.A(\add_x_19_5/n184 ));
   XOR2X4TS \add_x_19_5/U112  (.Y(\addr_calc/iir_write_addr[17] ), 
	.B(\add_x_19_5/n15 ), 
	.A(\add_x_19_5/n107 ));
   NAND2X1TS \add_x_19_5/U11  (.Y(\add_x_19_5/n37 ), 
	.B(FE_OFN559_offset_30_), 
	.A(FE_OFN239_addr_calc_iir_write_calc_count_30_));
   NAND2X1TS \add_x_19_5/U19  (.Y(\add_x_19_5/n42 ), 
	.B(FE_OFN347_offset_29_), 
	.A(n1851));
   NAND2X1TS \add_x_19_5/U29  (.Y(\add_x_19_5/n49 ), 
	.B(FE_OFN351_offset_28_), 
	.A(\addr_calc/iir_write_calc/count[28] ));
   NAND2X1TS \add_x_19_5/U39  (.Y(\add_x_19_5/n56 ), 
	.B(FE_OFN355_offset_27_), 
	.A(\addr_calc/iir_write_calc/count[27] ));
   NAND2X1TS \add_x_19_5/U45  (.Y(\add_x_19_5/n59 ), 
	.B(FE_OFN360_offset_26_), 
	.A(\addr_calc/iir_write_calc/count[26] ));
   NAND2X1TS \add_x_19_5/U53  (.Y(\add_x_19_5/n64 ), 
	.B(FE_OFN364_offset_25_), 
	.A(n1969));
   NAND2X2TS \add_x_19_5/U59  (.Y(\add_x_19_5/n67 ), 
	.B(FE_OFN367_offset_24_), 
	.A(n2051));
   NAND2X1TS \add_x_19_5/U74  (.Y(\add_x_19_5/n79 ), 
	.B(FE_OFN372_offset_23_), 
	.A(n1965));
   NAND2X6TS \add_x_19_5/U80  (.Y(\add_x_19_5/n82 ), 
	.B(FE_OCPUNCON1877_FE_OFN374_offset_22_), 
	.A(\addr_calc/iir_write_calc/count[22] ));
   NAND2X1TS \add_x_19_5/U88  (.Y(\add_x_19_5/n87 ), 
	.B(FE_OFN380_offset_21_), 
	.A(n1962));
   NAND2X1TS \add_x_19_5/U105  (.Y(\add_x_19_5/n98 ), 
	.B(FE_OFN384_offset_19_), 
	.A(n1958));
   NAND2X2TS \add_x_19_5/U111  (.Y(\add_x_19_5/n101 ), 
	.B(FE_OFN389_offset_18_), 
	.A(FE_OFN265_addr_calc_iir_write_calc_count_18_));
   NOR2X4TS \add_x_19_5/U52  (.Y(\add_x_19_5/n63 ), 
	.B(FE_OFN364_offset_25_), 
	.A(n1969));
   NOR2X4TS \add_x_19_5/U58  (.Y(\add_x_19_5/n66 ), 
	.B(FE_OFN367_offset_24_), 
	.A(n2051));
   NOR2X2TS \add_x_19_5/U87  (.Y(\add_x_19_5/n86 ), 
	.B(FE_OFN380_offset_21_), 
	.A(n1962));
   NOR2X2TS \add_x_19_5/U110  (.Y(\add_x_19_5/n100 ), 
	.B(FE_OFN389_offset_18_), 
	.A(FE_OFN265_addr_calc_iir_write_calc_count_18_));
   NOR2X8TS \add_x_19_5/U118  (.Y(\add_x_19_5/n105 ), 
	.B(FE_OFN392_offset_17_), 
	.A(\addr_calc/iir_write_calc/count[17] ));
   NOR2X2TS \add_x_19_5/U126  (.Y(\add_x_19_5/n110 ), 
	.B(FE_OFN397_offset_16_), 
	.A(\addr_calc/iir_write_calc/count[16] ));
   NAND2X1TS \add_x_19_5/U140  (.Y(\add_x_19_5/n121 ), 
	.B(FE_OCPUNCON1942_FE_OFN399_offset_15_), 
	.A(FE_OFN229_addr_calc_iir_write_calc_count_15_));
   NAND2X2TS \add_x_19_5/U146  (.Y(\add_x_19_5/n124 ), 
	.B(FE_OFN405_offset_14_), 
	.A(\addr_calc/iir_write_calc/count[14] ));
   NAND2X1TS \add_x_19_5/U154  (.Y(\add_x_19_5/n129 ), 
	.B(FE_OFN408_offset_13_), 
	.A(\addr_calc/iir_write_calc/count[13] ));
   NAND2X2TS \add_x_19_5/U160  (.Y(\add_x_19_5/n132 ), 
	.B(FE_OCPUNCON1073_FE_OFN410_offset_12_), 
	.A(\addr_calc/iir_write_calc/count[12] ));
   NAND2X2TS \add_x_19_5/U179  (.Y(\add_x_19_5/n145 ), 
	.B(FE_OFN421_offset_10_), 
	.A(\addr_calc/iir_write_calc/count[10] ));
   NAND2X2TS \add_x_19_5/U189  (.Y(\add_x_19_5/n152 ), 
	.B(FE_OFN424_offset_9_), 
	.A(\addr_calc/iir_write_calc/count[9] ));
   NAND2X8TS \add_x_19_5/U195  (.Y(\add_x_19_5/n155 ), 
	.B(\addr_calc/iir_write_calc/count[8] ), 
	.A(FE_OFN429_offset_8_));
   NOR2X4TS \add_x_19_5/U153  (.Y(\add_x_19_5/n128 ), 
	.B(FE_OFN408_offset_13_), 
	.A(\addr_calc/iir_write_calc/count[13] ));
   NOR2X2TS \add_x_19_5/U159  (.Y(\add_x_19_5/n131 ), 
	.B(FE_OCPUNCON1073_FE_OFN410_offset_12_), 
	.A(\addr_calc/iir_write_calc/count[12] ));
   NOR2X6TS \add_x_19_5/U178  (.Y(\add_x_19_5/n144 ), 
	.B(\addr_calc/iir_write_calc/count[10] ), 
	.A(FE_OFN421_offset_10_));
   NOR2X2TS \add_x_19_5/U194  (.Y(\add_x_19_5/n154 ), 
	.B(FE_OFN429_offset_8_), 
	.A(\addr_calc/iir_write_calc/count[8] ));
   NAND2X6TS \add_x_19_5/U206  (.Y(\add_x_19_5/n163 ), 
	.B(FE_OCP_RBN1840_offset_7_), 
	.A(n1683));
   NAND2X4TS \add_x_19_5/U228  (.Y(\add_x_19_5/n176 ), 
	.B(\addr_calc/iir_write_calc/count[4] ), 
	.A(FE_OFN444_offset_4_));
   NOR2X4TS \add_x_19_5/U211  (.Y(\add_x_19_5/n165 ), 
	.B(FE_OFN436_offset_6_), 
	.A(\addr_calc/iir_write_calc/count[6] ));
   NOR2X4TS \add_x_19_5/U227  (.Y(\add_x_19_5/n175 ), 
	.B(FE_OFN444_offset_4_), 
	.A(\addr_calc/iir_write_calc/count[4] ));
   NAND2X2TS \add_x_19_5/U237  (.Y(\add_x_19_5/n182 ), 
	.B(FE_OFN250_addr_calc_iir_write_calc_count_3_), 
	.A(FE_OCPUNCON1075_FE_OFN447_offset_3_));
   NAND2X8TS \add_x_19_5/U243  (.Y(\add_x_19_5/n185 ), 
	.B(\addr_calc/iir_write_calc/count[2] ), 
	.A(FE_OCPUNCON1076_FE_OFN451_offset_2_));
   NAND2X2TS \add_x_19_5/U250  (.Y(\add_x_19_5/n189 ), 
	.B(FE_OCP_RBN1919_offset_1_), 
	.A(\addr_calc/iir_write_calc/count[1] ));
   NOR2X8TS \add_x_19_5/U242  (.Y(\add_x_19_5/n184 ), 
	.B(FE_OCPUNCON1076_FE_OFN451_offset_2_), 
	.A(\addr_calc/iir_write_calc/count[2] ));
   NAND2X1TS \add_x_19_5/U247  (.Y(\add_x_19_5/n31 ), 
	.B(\add_x_19_5/n189 ), 
	.A(\add_x_19_5/n222 ));
   XNOR2X2TS \add_x_19_5/U229  (.Y(\addr_calc/iir_write_addr[3] ), 
	.B(\add_x_19_5/n29 ), 
	.A(\add_x_19_5/n183 ));
   NAND2X1TS \add_x_19_5/U234  (.Y(\add_x_19_5/n29 ), 
	.B(\add_x_19_5/n182 ), 
	.A(\add_x_19_5/n220 ));
   XNOR2X1TS \add_x_19_5/U221  (.Y(\addr_calc/iir_write_addr[4] ), 
	.B(\add_x_19_5/n28 ), 
	.A(n1818));
   NAND2X1TS \add_x_19_5/U225  (.Y(\add_x_19_5/n28 ), 
	.B(\add_x_19_5/n176 ), 
	.A(\add_x_19_5/n219 ));
   NAND2X1TS \add_x_19_5/U186  (.Y(\add_x_19_5/n23 ), 
	.B(\add_x_19_5/n152 ), 
	.A(\add_x_19_5/n214 ));
   NAND2X1TS \add_x_19_5/U176  (.Y(\add_x_19_5/n22 ), 
	.B(\add_x_19_5/n145 ), 
	.A(\add_x_19_5/n213 ));
   NAND2X2TS \add_x_19_5/U124  (.Y(\add_x_19_5/n16 ), 
	.B(\add_x_19_5/n111 ), 
	.A(\add_x_19_5/n207 ));
   XNOR2X4TS \add_x_19_5/U147  (.Y(\addr_calc/iir_write_addr[13] ), 
	.B(\add_x_19_5/n19 ), 
	.A(\add_x_19_5/n130 ));
   NAND2X1TS \add_x_19_5/U151  (.Y(\add_x_19_5/n19 ), 
	.B(\add_x_19_5/n129 ), 
	.A(\add_x_19_5/n210 ));
   NAND2X1TS \add_x_19_5/U116  (.Y(\add_x_19_5/n15 ), 
	.B(\add_x_19_5/n106 ), 
	.A(\add_x_19_5/n206 ));
   NAND2X1TS \add_x_19_5/U85  (.Y(\add_x_19_5/n11 ), 
	.B(\add_x_19_5/n87 ), 
	.A(\add_x_19_5/n202 ));
   NAND2X1TS \add_x_19_5/U26  (.Y(\add_x_19_5/n4 ), 
	.B(\add_x_19_5/n49 ), 
	.A(\add_x_19_5/n195 ));
   NAND2X1TS \add_x_19_5/U50  (.Y(\add_x_19_5/n7 ), 
	.B(\add_x_19_5/n64 ), 
	.A(\add_x_19_5/n198 ));
   NAND2X2TS \add_x_19_5/U119  (.Y(\add_x_19_5/n106 ), 
	.B(FE_OFN392_offset_17_), 
	.A(\addr_calc/iir_write_calc/count[17] ));
   NAND2X1TS \add_x_19_5/U32  (.Y(\add_x_19_5/n51 ), 
	.B(\add_x_19_5/n53 ), 
	.A(\add_x_19_5/n61 ));
   NAND2X4TS \add_x_19_5/U98  (.Y(\add_x_19_5/n93 ), 
	.B(\add_x_19_5/n95 ), 
	.A(\add_x_19_5/n103 ));
   NAND2X1TS \add_x_19_5/U171  (.Y(\add_x_19_5/n140 ), 
	.B(FE_OFN417_offset_11_), 
	.A(\addr_calc/iir_write_calc/count[11] ));
   NAND2X4TS \add_x_19_5/U164  (.Y(\add_x_19_5/n135 ), 
	.B(\add_x_19_5/n137 ), 
	.A(\add_x_19_5/n149 ));
   NAND2X4TS \add_x_19_5/U220  (.Y(\add_x_19_5/n171 ), 
	.B(n1686), 
	.A(FE_OCP_RBN1492_offset_5_));
   NOR2X4TS \add_x_19_0/U219  (.Y(\add_x_19_0/n170 ), 
	.B(FE_OCP_RBN1495_offset_5_), 
	.A(FE_OFN251_addr_calc_fft_read_calc_count_5_));
   NAND2X6TS \add_x_19_0/U127  (.Y(\add_x_19_0/n111 ), 
	.B(FE_OFN396_offset_16_), 
	.A(\addr_calc/fft_read_calc/count[16] ));
   AOI21X1TS \add_x_19_0/U214  (.Y(\add_x_19_0/n167 ), 
	.B0(\add_x_19_0/n169 ), 
	.A1(\add_x_19_0/n168 ), 
	.A0(\add_x_19_0/n177 ));
   XOR2X1TS \add_x_19_0/U190  (.Y(\addr_calc/fft_read_addr[8] ), 
	.B(\add_x_19_0/n24 ), 
	.A(\add_x_19_0/n156 ));
   OAI21X1TS \add_x_19_0/U142  (.Y(\add_x_19_0/n122 ), 
	.B0(\add_x_19_0/n124 ), 
	.A1(\add_x_19_0/n123 ), 
	.A0(\add_x_19_0/n125 ));
   AOI21X4TS \add_x_19_0/U113  (.Y(\add_x_19_0/n102 ), 
	.B0(\add_x_19_0/n104 ), 
	.A1(\add_x_19_0/n103 ), 
	.A0(\add_x_19_0/n112 ));
   OAI21X4TS \add_x_19_0/U31  (.Y(\add_x_19_0/n50 ), 
	.B0(\add_x_19_0/n52 ), 
	.A1(\add_x_19_0/n51 ), 
	.A0(\add_x_19_0/n68 ));
   NOR2X1TS \add_x_19_0/U10  (.Y(\add_x_19_0/n36 ), 
	.B(FE_OFN344_offset_30_), 
	.A(FE_OFN278_addr_calc_fft_read_calc_count_30_));
   AOI21X4TS \add_x_19_0/U23  (.Y(\add_x_19_0/n45 ), 
	.B0(\add_x_19_0/n47 ), 
	.A1(\add_x_19_0/n46 ), 
	.A0(\add_x_19_0/n73 ));
   OAI21X2TS \add_x_19_0/U25  (.Y(\add_x_19_0/n47 ), 
	.B0(\add_x_19_0/n49 ), 
	.A1(\add_x_19_0/n48 ), 
	.A0(\add_x_19_0/n52 ));
   OAI21X1TS \add_x_19_0/U35  (.Y(\add_x_19_0/n54 ), 
	.B0(\add_x_19_0/n56 ), 
	.A1(\add_x_19_0/n59 ), 
	.A0(\add_x_19_0/n55 ));
   OAI21X2TS \add_x_19_0/U49  (.Y(\add_x_19_0/n62 ), 
	.B0(\add_x_19_0/n64 ), 
	.A1(\add_x_19_0/n67 ), 
	.A0(\add_x_19_0/n63 ));
   OAI21X4TS \add_x_19_0/U115  (.Y(\add_x_19_0/n104 ), 
	.B0(\add_x_19_0/n106 ), 
	.A1(\add_x_19_0/n111 ), 
	.A0(\add_x_19_0/n105 ));
   NOR2X4TS \add_x_19_0/U69  (.Y(\add_x_19_0/n76 ), 
	.B(\add_x_19_0/n78 ), 
	.A(\add_x_19_0/n81 ));
   NOR2X2TS \add_x_19_0/U100  (.Y(\add_x_19_0/n95 ), 
	.B(\add_x_19_0/n97 ), 
	.A(\add_x_19_0/n100 ));
   NOR2X2TS \add_x_19_0/U114  (.Y(\add_x_19_0/n103 ), 
	.B(\add_x_19_0/n105 ), 
	.A(\add_x_19_0/n110 ));
   OAI21X2TS \add_x_19_0/U185  (.Y(\add_x_19_0/n150 ), 
	.B0(\add_x_19_0/n152 ), 
	.A1(\add_x_19_0/n155 ), 
	.A0(\add_x_19_0/n151 ));
   NOR2X2TS \add_x_19_0/U166  (.Y(\add_x_19_0/n137 ), 
	.B(\add_x_19_0/n139 ), 
	.A(\add_x_19_0/n144 ));
   NOR2X4TS \add_x_19_0/U170  (.Y(\add_x_19_0/n139 ), 
	.B(\addr_calc/fft_read_calc/count[11] ), 
	.A(FE_OCPUNCON656_FE_OFN414_offset_11_));
   NOR2X1TS \add_x_19_0/U184  (.Y(\add_x_19_0/n149 ), 
	.B(\add_x_19_0/n154 ), 
	.A(\add_x_19_0/n151 ));
   OAI21X4TS \add_x_19_0/U216  (.Y(\add_x_19_0/n169 ), 
	.B0(\add_x_19_0/n171 ), 
	.A1(\add_x_19_0/n170 ), 
	.A0(\add_x_19_0/n176 ));
   NOR2X4TS \add_x_19_0/U215  (.Y(\add_x_19_0/n168 ), 
	.B(\add_x_19_0/n170 ), 
	.A(\add_x_19_0/n175 ));
   XOR2X4TS \add_x_19_0/U112  (.Y(\addr_calc/fft_read_addr[17] ), 
	.B(\add_x_19_0/n15 ), 
	.A(\add_x_19_0/n107 ));
   NAND2X1TS \add_x_19_0/U11  (.Y(\add_x_19_0/n37 ), 
	.B(FE_OFN344_offset_30_), 
	.A(FE_OFN278_addr_calc_fft_read_calc_count_30_));
   NAND2X1TS \add_x_19_0/U19  (.Y(\add_x_19_0/n42 ), 
	.B(FE_OFN348_offset_29_), 
	.A(FE_OFN275_addr_calc_fft_read_calc_count_29_));
   NAND2X1TS \add_x_19_0/U29  (.Y(\add_x_19_0/n49 ), 
	.B(FE_OFN352_offset_28_), 
	.A(n2559));
   NAND2X1TS \add_x_19_0/U39  (.Y(\add_x_19_0/n56 ), 
	.B(FE_OFN356_offset_27_), 
	.A(n1944));
   NAND2X1TS \add_x_19_0/U45  (.Y(\add_x_19_0/n59 ), 
	.B(FE_OFN359_offset_26_), 
	.A(\addr_calc/fft_read_calc/count[26] ));
   NAND2X1TS \add_x_19_0/U53  (.Y(\add_x_19_0/n64 ), 
	.B(FE_OFN363_offset_25_), 
	.A(n1947));
   NAND2X2TS \add_x_19_0/U59  (.Y(\add_x_19_0/n67 ), 
	.B(FE_OFN368_offset_24_), 
	.A(n2038));
   NAND2X1TS \add_x_19_0/U74  (.Y(\add_x_19_0/n79 ), 
	.B(FE_OFN371_offset_23_), 
	.A(n1950));
   NAND2X2TS \add_x_19_0/U80  (.Y(\add_x_19_0/n82 ), 
	.B(FE_OFN375_offset_22_), 
	.A(\addr_calc/fft_read_calc/count[22] ));
   NAND2X1TS \add_x_19_0/U88  (.Y(\add_x_19_0/n87 ), 
	.B(FE_OCPUNCON1078_FE_OFN377_offset_21_), 
	.A(FE_OFN288_addr_calc_fft_read_calc_count_21_));
   NAND2X1TS \add_x_19_0/U105  (.Y(\add_x_19_0/n98 ), 
	.B(FE_OCPUNCON1079_FE_OFN382_offset_19_), 
	.A(n1956));
   NAND2X2TS \add_x_19_0/U111  (.Y(\add_x_19_0/n101 ), 
	.B(FE_OCPUNCON1080_FE_OFN386_offset_18_), 
	.A(\addr_calc/fft_read_calc/count[18] ));
   NAND2X1TS \add_x_19_0/U119  (.Y(\add_x_19_0/n106 ), 
	.B(FE_OFN393_offset_17_), 
	.A(FE_OFN287_addr_calc_fft_read_calc_count_17_));
   NOR2X4TS \add_x_19_0/U52  (.Y(\add_x_19_0/n63 ), 
	.B(FE_OFN363_offset_25_), 
	.A(n1947));
   NOR2X2TS \add_x_19_0/U79  (.Y(\add_x_19_0/n81 ), 
	.B(FE_OFN375_offset_22_), 
	.A(n1665));
   NOR2X4TS \add_x_19_0/U87  (.Y(\add_x_19_0/n86 ), 
	.B(FE_OCPUNCON1078_FE_OFN377_offset_21_), 
	.A(FE_OFN288_addr_calc_fft_read_calc_count_21_));
   NOR2X2TS \add_x_19_0/U110  (.Y(\add_x_19_0/n100 ), 
	.B(\addr_calc/fft_read_calc/count[18] ), 
	.A(FE_OCPUNCON1080_FE_OFN386_offset_18_));
   NOR2X8TS \add_x_19_0/U118  (.Y(\add_x_19_0/n105 ), 
	.B(FE_OFN287_addr_calc_fft_read_calc_count_17_), 
	.A(FE_OFN393_offset_17_));
   NAND2X1TS \add_x_19_0/U140  (.Y(\add_x_19_0/n121 ), 
	.B(FE_OFN400_offset_15_), 
	.A(n1689));
   NAND2X1TS \add_x_19_0/U146  (.Y(\add_x_19_0/n124 ), 
	.B(FE_OFN404_offset_14_), 
	.A(n2043));
   NAND2X1TS \add_x_19_0/U154  (.Y(\add_x_19_0/n129 ), 
	.B(FE_OCPUNCON1943_FE_OFN407_offset_13_), 
	.A(n1967));
   NAND2X2TS \add_x_19_0/U179  (.Y(\add_x_19_0/n145 ), 
	.B(\addr_calc/fft_read_calc/count[10] ), 
	.A(FE_OCPUNCON657_FE_OFN418_offset_10_));
   NAND2X1TS \add_x_19_0/U189  (.Y(\add_x_19_0/n152 ), 
	.B(\addr_calc/fft_read_calc/count[9] ), 
	.A(FE_OCPUNCON658_FE_OFN422_offset_9_));
   NAND2X2TS \add_x_19_0/U195  (.Y(\add_x_19_0/n155 ), 
	.B(\addr_calc/fft_read_calc/count[8] ), 
	.A(FE_OFN428_offset_8_));
   NOR2X4TS \add_x_19_0/U188  (.Y(\add_x_19_0/n151 ), 
	.B(FE_OCPUNCON658_FE_OFN422_offset_9_), 
	.A(\addr_calc/fft_read_calc/count[9] ));
   NOR2X1TS \add_x_19_0/U194  (.Y(\add_x_19_0/n154 ), 
	.B(\addr_calc/fft_read_calc/count[8] ), 
	.A(FE_OFN428_offset_8_));
   NAND2X2TS \add_x_19_0/U206  (.Y(\add_x_19_0/n163 ), 
	.B(n1666), 
	.A(FE_OCPUNCON1278_offset_7_));
   NAND2X1TS \add_x_19_0/U212  (.Y(\add_x_19_0/n166 ), 
	.B(FE_OCPUNCON726_FE_OFN435_offset_6_), 
	.A(FE_OFN225_addr_calc_fft_read_calc_count_6_));
   NAND2X2TS \add_x_19_0/U228  (.Y(\add_x_19_0/n176 ), 
	.B(FE_OFN264_addr_calc_fft_read_calc_count_4_), 
	.A(FE_OCPUNCON1425_FE_OFN443_offset_4_));
   NAND2X4TS \add_x_19_0/U237  (.Y(\add_x_19_0/n182 ), 
	.B(FE_OFN449_offset_3_), 
	.A(\addr_calc/fft_read_calc/count[3] ));
   NAND2X4TS \add_x_19_0/U243  (.Y(\add_x_19_0/n185 ), 
	.B(FE_OFN452_offset_2_), 
	.A(\addr_calc/fft_read_calc/count[2] ));
   NAND2X2TS \add_x_19_0/U250  (.Y(\add_x_19_0/n189 ), 
	.B(FE_OCPUNCON1874_offset_1_), 
	.A(\addr_calc/fft_read_calc/count[1] ));
   XNOR2X1TS \add_x_19_0/U221  (.Y(\addr_calc/fft_read_addr[4] ), 
	.B(\add_x_19_0/n28 ), 
	.A(\add_x_19_0/n177 ));
   NAND2X1TS \add_x_19_0/U225  (.Y(\add_x_19_0/n28 ), 
	.B(\add_x_19_0/n176 ), 
	.A(\add_x_19_0/n219 ));
   NAND2X1TS \add_x_19_0/U192  (.Y(\add_x_19_0/n24 ), 
	.B(\add_x_19_0/n155 ), 
	.A(\add_x_19_0/n215 ));
   XNOR2XLTS \add_x_19_0/U172  (.Y(\addr_calc/fft_read_addr[10] ), 
	.B(\add_x_19_0/n22 ), 
	.A(\add_x_19_0/n146 ));
   NAND2X1TS \add_x_19_0/U176  (.Y(\add_x_19_0/n22 ), 
	.B(\add_x_19_0/n145 ), 
	.A(\add_x_19_0/n213 ));
   XNOR2X4TS \add_x_19_0/U147  (.Y(\addr_calc/fft_read_addr[13] ), 
	.B(\add_x_19_0/n19 ), 
	.A(\add_x_19_0/n130 ));
   NAND2X1TS \add_x_19_0/U151  (.Y(\add_x_19_0/n19 ), 
	.B(\add_x_19_0/n129 ), 
	.A(\add_x_19_0/n210 ));
   XNOR2X2TS \add_x_19_0/U128  (.Y(\addr_calc/fft_read_addr[15] ), 
	.B(\add_x_19_0/n17 ), 
	.A(\add_x_19_0/n122 ));
   NAND2X1TS \add_x_19_0/U137  (.Y(\add_x_19_0/n17 ), 
	.B(\add_x_19_0/n121 ), 
	.A(\add_x_19_0/n208 ));
   NAND2X1TS \add_x_19_0/U116  (.Y(\add_x_19_0/n15 ), 
	.B(\add_x_19_0/n106 ), 
	.A(\add_x_19_0/n206 ));
   XNOR2X4TS \add_x_19_0/U95  (.Y(\addr_calc/fft_read_addr[19] ), 
	.B(\add_x_19_0/n13 ), 
	.A(\add_x_19_0/n99 ));
   NAND2X1TS \add_x_19_0/U102  (.Y(\add_x_19_0/n13 ), 
	.B(\add_x_19_0/n98 ), 
	.A(\add_x_19_0/n204 ));
   NAND2X1TS \add_x_19_0/U85  (.Y(\add_x_19_0/n11 ), 
	.B(\add_x_19_0/n87 ), 
	.A(\add_x_19_0/n202 ));
   NAND2X2TS \add_x_19_0/U26  (.Y(\add_x_19_0/n4 ), 
	.B(\add_x_19_0/n49 ), 
	.A(\add_x_19_0/n195 ));
   XNOR2X4TS \add_x_19_0/U46  (.Y(\addr_calc/fft_read_addr[25] ), 
	.B(\add_x_19_0/n7 ), 
	.A(\add_x_19_0/n65 ));
   NAND2X1TS \add_x_19_0/U50  (.Y(\add_x_19_0/n7 ), 
	.B(\add_x_19_0/n64 ), 
	.A(\add_x_19_0/n198 ));
   NAND2X4TS \add_x_19_0/U2  (.Y(\add_x_19_0/n1 ), 
	.B(\add_x_19_0/n34 ), 
	.A(n2627));
   NAND2X4TS \add_x_19_0/U22  (.Y(\add_x_19_0/n44 ), 
	.B(\add_x_19_0/n72 ), 
	.A(\add_x_19_0/n46 ));
   NAND2X2TS \add_x_19_0/U32  (.Y(\add_x_19_0/n51 ), 
	.B(\add_x_19_0/n53 ), 
	.A(\add_x_19_0/n61 ));
   NAND2X4TS \add_x_19_0/U98  (.Y(\add_x_19_0/n93 ), 
	.B(\add_x_19_0/n95 ), 
	.A(\add_x_19_0/n103 ));
   NAND2X1TS \add_x_19_0/U171  (.Y(\add_x_19_0/n140 ), 
	.B(FE_OCPUNCON656_FE_OFN414_offset_11_), 
	.A(\addr_calc/fft_read_calc/count[11] ));
   NAND2X4TS \add_x_19_0/U164  (.Y(\add_x_19_0/n135 ), 
	.B(\add_x_19_0/n137 ), 
	.A(\add_x_19_0/n149 ));
   NAND2X1TS \add_x_19_0/U220  (.Y(\add_x_19_0/n171 ), 
	.B(FE_OCP_RBN1495_offset_5_), 
	.A(FE_OFN251_addr_calc_fft_read_calc_count_5_));
   NOR2X1TS \DP_OP_159_297_3515/U1098  (.Y(\DP_OP_159_297_3515/n1051 ), 
	.B(\DP_OP_159_297_3515/n1052 ), 
	.A(\DP_OP_159_297_3515/n1063 ));
   NAND2X1TS \DP_OP_159_297_3515/U964  (.Y(\DP_OP_159_297_3515/n959 ), 
	.B(FE_OFN477_filesize_20_), 
	.A(FE_OFN478_filesize_19_));
   NOR2XLTS \DP_OP_159_297_3515/U1050  (.Y(\DP_OP_159_297_3515/n1018 ), 
	.B(\DP_OP_159_297_3515/n873 ), 
	.A(\DP_OP_159_297_3515/n1026 ));
   NAND2X1TS \DP_OP_159_297_3515/U990  (.Y(\DP_OP_159_297_3515/n976 ), 
	.B(n2369), 
	.A(FE_OFN553_n1789));
   NOR2X1TS \DP_OP_159_297_3515/U798  (.Y(\DP_OP_159_297_3515/n764 ), 
	.B(\DP_OP_159_297_3515/n766 ), 
	.A(\DP_OP_159_297_3515/n768 ));
   NOR2X1TS \DP_OP_159_297_3515/U810  (.Y(\DP_OP_159_297_3515/n774 ), 
	.B(\DP_OP_159_297_3515/n778 ), 
	.A(\DP_OP_159_297_3515/n776 ));
   NOR2X1TS \DP_OP_159_297_3515/U757  (.Y(\DP_OP_159_297_3515/n728 ), 
	.B(\DP_OP_159_297_3515/n737 ), 
	.A(\DP_OP_159_297_3515/n730 ));
   NOR2X1TS \DP_OP_159_297_3515/U1030  (.Y(\DP_OP_159_297_3515/n1004 ), 
	.B(\DP_OP_159_297_3515/n871 ), 
	.A(\DP_OP_159_297_3515/n1012 ));
   NOR2X1TS \DP_OP_159_297_3515/U1020  (.Y(\DP_OP_159_297_3515/n997 ), 
	.B(\DP_OP_159_297_3515/n998 ), 
	.A(\DP_OP_159_297_3515/n1012 ));
   NOR2X1TS \DP_OP_159_297_3515/U971  (.Y(\DP_OP_159_297_3515/n963 ), 
	.B(\DP_OP_159_297_3515/n964 ), 
	.A(\DP_OP_159_297_3515/n971 ));
   NOR2X1TS \DP_OP_159_297_3515/U861  (.Y(\DP_OP_159_297_3515/n886 ), 
	.B(\DP_OP_159_297_3515/n887 ), 
	.A(FE_OFN114_DP_OP_159_297_3515_n852));
   NOR2X1TS \DP_OP_159_297_3515/U871  (.Y(\DP_OP_159_297_3515/n893 ), 
	.B(\DP_OP_159_297_3515/n894 ), 
	.A(FE_OFN114_DP_OP_159_297_3515_n852));
   NOR2X1TS \DP_OP_159_297_3515/U931  (.Y(\DP_OP_159_297_3515/n935 ), 
	.B(\DP_OP_159_297_3515/n936 ), 
	.A(\DP_OP_159_297_3515/n957 ));
   NOR2X1TS \DP_OP_159_297_3515/U951  (.Y(\DP_OP_159_297_3515/n949 ), 
	.B(\DP_OP_159_297_3515/n950 ), 
	.A(\DP_OP_159_297_3515/n957 ));
   NOR2X1TS \DP_OP_159_297_3515/U891  (.Y(\DP_OP_159_297_3515/n907 ), 
	.B(\DP_OP_159_297_3515/n908 ), 
	.A(FE_OFN114_DP_OP_159_297_3515_n852));
   NOR2X1TS \DP_OP_159_297_3515/U901  (.Y(\DP_OP_159_297_3515/n914 ), 
	.B(\DP_OP_159_297_3515/n915 ), 
	.A(\DP_OP_159_297_3515/n852 ));
   NAND2X1TS \DP_OP_159_297_3515/U791  (.Y(\DP_OP_159_297_3515/n758 ), 
	.B(n2606), 
	.A(\DP_OP_159_297_3515/n764 ));
   XNOR2X1TS \DP_OP_159_297_3515/U800  (.Y(\DP_OP_159_297_3515/n766 ), 
	.B(FE_OFN250_addr_calc_iir_write_calc_count_3_), 
	.A(n2611));
   NAND2X1TS \DP_OP_159_297_3515/U803  (.Y(\DP_OP_159_297_3515/n768 ), 
	.B(n2604), 
	.A(\DP_OP_159_297_3515/n774 ));
   XNOR2X1TS \DP_OP_159_297_3515/U812  (.Y(\DP_OP_159_297_3515/n776 ), 
	.B(\addr_calc/iir_write_calc/count[1] ), 
	.A(FE_OFN501_filesize_1_));
   NAND2X1TS \DP_OP_159_297_3515/U773  (.Y(\DP_OP_159_297_3515/n742 ), 
	.B(n2626), 
	.A(n2605));
   XNOR2X1TS \DP_OP_159_297_3515/U767  (.Y(\DP_OP_159_297_3515/n737 ), 
	.B(\addr_calc/iir_write_calc/count[7] ), 
	.A(n2609));
   NAND2X1TS \DP_OP_159_297_3515/U1088  (.Y(\DP_OP_159_297_3515/n1044 ), 
	.B(n2362), 
	.A(\DP_OP_159_297_3515/n1051 ));
   NAND2X1TS \DP_OP_159_297_3515/U1011  (.Y(\DP_OP_159_297_3515/n991 ), 
	.B(FE_OFN484_filesize_15_), 
	.A(\DP_OP_159_297_3515/n999 ));
   NAND2X1TS \DP_OP_159_297_3515/U860  (.Y(\DP_OP_159_297_3515/n885 ), 
	.B(\DP_OP_159_297_3515/n886 ), 
	.A(FE_OCPUNCON1566_n1789));
   NAND2X1TS \DP_OP_159_297_3515/U862  (.Y(\DP_OP_159_297_3515/n887 ), 
	.B(n2603), 
	.A(\DP_OP_159_297_3515/n902 ));
   NAND2X1TS \DP_OP_159_297_3515/U872  (.Y(\DP_OP_159_297_3515/n894 ), 
	.B(FE_OFN465_filesize_29_), 
	.A(\DP_OP_159_297_3515/n902 ));
   NAND2X1TS \DP_OP_159_297_3515/U932  (.Y(\DP_OP_159_297_3515/n936 ), 
	.B(FE_OFN473_filesize_23_), 
	.A(\DP_OP_159_297_3515/n944 ));
   NAND2X1TS \DP_OP_159_297_3515/U892  (.Y(\DP_OP_159_297_3515/n908 ), 
	.B(FE_OFN467_filesize_27_), 
	.A(\DP_OP_159_297_3515/n916 ));
   NAND2X1TS \DP_OP_159_297_3515/U924  (.Y(\DP_OP_159_297_3515/n931 ), 
	.B(FE_OFN471_filesize_24_), 
	.A(FE_OFN472_filesize_23_));
   NOR2X2TS \DP_OP_158_296_6262/U305  (.Y(\DP_OP_158_296_6262/n280 ), 
	.B(FE_OFN539_DP_OP_158_296_6262_n318), 
	.A(\DP_OP_158_296_6262/n282 ));
   NOR2X1TS \DP_OP_158_296_6262/U379  (.Y(\DP_OP_158_296_6262/n347 ), 
	.B(\DP_OP_158_296_6262/n365 ), 
	.A(\DP_OP_158_296_6262/n349 ));
   NOR2X1TS \DP_OP_158_296_6262/U406  (.Y(\DP_OP_158_296_6262/n371 ), 
	.B(\DP_OP_158_296_6262/n375 ), 
	.A(\DP_OP_158_296_6262/n373 ));
   NOR2X1TS \DP_OP_158_296_6262/U309  (.Y(\DP_OP_158_296_6262/n284 ), 
	.B(\DP_OP_158_296_6262/n286 ), 
	.A(\DP_OP_158_296_6262/n297 ));
   NOR2X1TS \DP_OP_158_296_6262/U1803  (.Y(\DP_OP_158_296_6262/n1828 ), 
	.B(\DP_OP_158_296_6262/n1829 ), 
	.A(\DP_OP_158_296_6262/n1792 ));
   NAND2X1TS \DP_OP_158_296_6262/U399  (.Y(\DP_OP_158_296_6262/n365 ), 
	.B(n2590), 
	.A(\DP_OP_158_296_6262/n371 ));
   XNOR2X1TS \DP_OP_158_296_6262/U408  (.Y(\DP_OP_158_296_6262/n373 ), 
	.B(FE_OFN249_addr_calc_fir_read_calc_count_1_), 
	.A(n2597));
   NAND2X1TS \DP_OP_158_296_6262/U381  (.Y(\DP_OP_158_296_6262/n349 ), 
	.B(n2600), 
	.A(n2592));
   NAND2X1TS \DP_OP_158_296_6262/U359  (.Y(\DP_OP_158_296_6262/n329 ), 
	.B(n2591), 
	.A(n2601));
   XNOR2X1TS \DP_OP_158_296_6262/U351  (.Y(\DP_OP_158_296_6262/n322 ), 
	.B(FE_OFN227_addr_calc_fir_read_calc_count_7_), 
	.A(n1651));
   NAND2X1TS \DP_OP_158_296_6262/U307  (.Y(\DP_OP_158_296_6262/n282 ), 
	.B(\DP_OP_158_296_6262/n304 ), 
	.A(\DP_OP_158_296_6262/n284 ));
   XNOR2X1TS \DP_OP_158_296_6262/U343  (.Y(\DP_OP_158_296_6262/n315 ), 
	.B(n1997), 
	.A(n2598));
   XNOR2X1TS \DP_OP_158_296_6262/U333  (.Y(\DP_OP_158_296_6262/n306 ), 
	.B(n1900), 
	.A(n1469));
   XNOR2X1TS \DP_OP_158_296_6262/U311  (.Y(\DP_OP_158_296_6262/n286 ), 
	.B(n1895), 
	.A(n1660));
   XNOR2X1TS \DP_OP_158_296_6262/U263  (.Y(\DP_OP_158_296_6262/n242 ), 
	.B(n1890), 
	.A(n1658));
   XNOR2X1TS \DP_OP_158_296_6262/U277  (.Y(\DP_OP_158_296_6262/n255 ), 
	.B(n1690), 
	.A(n1657));
   XNOR2X1TS \DP_OP_158_296_6262/U289  (.Y(\DP_OP_158_296_6262/n266 ), 
	.B(n1893), 
	.A(FE_OFN524_n1659));
   XNOR2X1TS \DP_OP_158_296_6262/U250  (.Y(\DP_OP_158_296_6262/n230 ), 
	.B(n1888), 
	.A(n2594));
   XNOR2X1TS \DP_OP_158_296_6262/U10  (.Y(\DP_OP_158_296_6262/n5 ), 
	.B(\addr_calc/fir_read_calc/count[31] ), 
	.A(n1778));
   NAND2X1TS \DP_OP_158_296_6262/U2032  (.Y(\DP_OP_158_296_6262/n2004 ), 
	.B(\DP_OP_159_297_3515/n880 ), 
	.A(\DP_OP_158_296_6262/n2010 ));
   NAND2X1TS \DP_OP_158_296_6262/U1981  (.Y(\DP_OP_158_296_6262/n1965 ), 
	.B(\DP_OP_158_296_6262/n1966 ), 
	.A(n1138));
   NAND2X1TS \DP_OP_158_296_6262/U1945  (.Y(\DP_OP_158_296_6262/n1937 ), 
	.B(\DP_OP_158_296_6262/n1959 ), 
	.A(\DP_OP_158_296_6262/n1938 ));
   NAND2XLTS \DP_OP_158_296_6262/U1963  (.Y(\DP_OP_158_296_6262/n1951 ), 
	.B(\DP_OP_158_296_6262/n1952 ), 
	.A(\DP_OP_158_296_6262/n1959 ));
   NAND2X1TS \DP_OP_158_296_6262/U1910  (.Y(\DP_OP_158_296_6262/n1910 ), 
	.B(\DP_OP_158_296_6262/n1911 ), 
	.A(\DP_OP_158_296_6262/n1918 ));
   NAND2X1TS \DP_OP_158_296_6262/U1802  (.Y(\DP_OP_158_296_6262/n1827 ), 
	.B(\DP_OP_158_296_6262/n1828 ), 
	.A(FE_OFN113_DP_OP_158_296_6262_n1791));
   NAND2X1TS \DP_OP_158_296_6262/U1838  (.Y(\DP_OP_158_296_6262/n1854 ), 
	.B(FE_OFN112_DP_OP_158_296_6262_n1791), 
	.A(\DP_OP_158_296_6262/n1855 ));
   NAND2XLTS \DP_OP_158_296_6262/U1892  (.Y(\DP_OP_158_296_6262/n1896 ), 
	.B(\DP_OP_158_296_6262/n1897 ), 
	.A(\DP_OP_158_296_6262/n1904 ));
   NOR2X1TS \add_x_22_4/U101  (.Y(\add_x_22_4/n81 ), 
	.B(\add_x_22_4/n84 ), 
	.A(\add_x_22_4/n85 ));
   NOR2X1TS \add_x_22_4/U127  (.Y(\add_x_22_4/n102 ), 
	.B(\add_x_22_4/n103 ), 
	.A(\add_x_22_4/n110 ));
   NOR2X1TS \add_x_22_4/U132  (.Y(\add_x_22_4/n106 ), 
	.B(\add_x_22_4/n109 ), 
	.A(\add_x_22_4/n110 ));
   NOR2X1TS \add_x_22_4/U85  (.Y(\add_x_22_4/n68 ), 
	.B(\add_x_22_4/n69 ), 
	.A(\add_x_22_4/n76 ));
   NOR2X1TS \add_x_22_4/U63  (.Y(\add_x_22_4/n50 ), 
	.B(\add_x_22_4/n51 ), 
	.A(\add_x_22_4/n58 ));
   NOR2X1TS \add_x_22_4/U21  (.Y(\add_x_22_4/n16 ), 
	.B(\add_x_22_4/n17 ), 
	.A(\add_x_22_4/n24 ));
   NOR2X1TS \add_x_22_4/U12  (.Y(\add_x_22_4/n9 ), 
	.B(\add_x_22_4/n10 ), 
	.A(\add_x_22_4/n17 ));
   NOR2X1TS \add_x_22_4/U34  (.Y(\add_x_22_4/n27 ), 
	.B(\add_x_22_4/n28 ), 
	.A(\add_x_22_4/n35 ));
   NOR2X1TS \add_x_22_4/U68  (.Y(\add_x_22_4/n54 ), 
	.B(\add_x_22_4/n57 ), 
	.A(\add_x_22_4/n58 ));
   NOR2X1TS \add_x_22_4/U43  (.Y(\add_x_22_4/n34 ), 
	.B(\add_x_22_4/n35 ), 
	.A(\add_x_22_4/n42 ));
   NOR2X1TS \add_x_22_4/U54  (.Y(\add_x_22_4/n43 ), 
	.B(\add_x_22_4/n44 ), 
	.A(\add_x_22_4/n51 ));
   NOR2X1TS \add_x_22_4/U138  (.Y(\add_x_22_4/n111 ), 
	.B(\add_x_22_4/n119 ), 
	.A(\add_x_22_4/n112 ));
   NOR2X1TS \add_x_22_4/U96  (.Y(\add_x_22_4/n77 ), 
	.B(\add_x_22_4/n78 ), 
	.A(\add_x_22_4/n87 ));
   XNOR2X1TS \add_x_22_4/U142  (.Y(\addr_calc/iir_read_calc/counter/N45 ), 
	.B(\add_x_22_4/n117 ), 
	.A(\add_x_22_4/n118 ));
   XNOR2X1TS \add_x_22_4/U146  (.Y(\addr_calc/iir_read_calc/counter/N44 ), 
	.B(n2580), 
	.A(\add_x_22_4/n121 ));
   XNOR2X1TS \add_x_22_4/U80  (.Y(\addr_calc/iir_read_calc/counter/N57 ), 
	.B(\add_x_22_4/n67 ), 
	.A(\add_x_22_4/n68 ));
   NAND2X1TS \add_x_22_4/U143  (.Y(\add_x_22_4/n115 ), 
	.B(n2015), 
	.A(\add_x_22_4/n118 ));
   XNOR2X1TS \add_x_22_4/U58  (.Y(\addr_calc/iir_read_calc/counter/N61 ), 
	.B(n2024), 
	.A(\add_x_22_4/n50 ));
   XNOR2X1TS \add_x_22_4/U47  (.Y(\addr_calc/iir_read_calc/counter/N63 ), 
	.B(n2027), 
	.A(\add_x_22_4/n41 ));
   XNOR2X1TS \add_x_22_4/U89  (.Y(\addr_calc/iir_read_calc/counter/N55 ), 
	.B(\add_x_22_4/n74 ), 
	.A(\add_x_22_4/n75 ));
   XNOR2X1TS \add_x_22_4/U93  (.Y(\addr_calc/iir_read_calc/counter/N54 ), 
	.B(\add_x_22_4/n80 ), 
	.A(\add_x_22_4/n81 ));
   NAND2X1TS \add_x_22_4/U123  (.Y(\add_x_22_4/n99 ), 
	.B(n2018), 
	.A(\add_x_22_4/n102 ));
   XNOR2X1TS \add_x_22_4/U126  (.Y(\addr_calc/iir_read_calc/counter/N48 ), 
	.B(\add_x_22_4/n105 ), 
	.A(\add_x_22_4/n106 ));
   XNOR2X1TS \add_x_22_4/U111  (.Y(\addr_calc/iir_read_calc/counter/N51 ), 
	.B(\add_x_22_4/n92 ), 
	.A(\add_x_22_4/n93 ));
   NAND2X1TS \add_x_22_4/U81  (.Y(\add_x_22_4/n65 ), 
	.B(n1784), 
	.A(\add_x_22_4/n68 ));
   NAND2X1TS \add_x_22_4/U95  (.Y(\add_x_22_4/n76 ), 
	.B(\add_x_22_4/n77 ), 
	.A(\add_x_22_4/n93 ));
   NAND2X1TS \add_x_22_4/U11  (.Y(\add_x_22_4/n8 ), 
	.B(\add_x_22_4/n9 ), 
	.A(\add_x_22_4/n23 ));
   NAND2X1TS \add_x_22_4/U59  (.Y(\add_x_22_4/n47 ), 
	.B(\addr_calc/iir_read_calc/count[18] ), 
	.A(\add_x_22_4/n50 ));
   NAND2X1TS \add_x_22_4/U26  (.Y(\add_x_22_4/n20 ), 
	.B(n2034), 
	.A(\add_x_22_4/n23 ));
   XNOR2X1TS \add_x_22_4/U25  (.Y(\addr_calc/iir_read_calc/counter/N67 ), 
	.B(n2033), 
	.A(\add_x_22_4/n23 ));
   ADDHXLTS \add_x_22_4/U2  (.S(\addr_calc/iir_read_calc/counter/N73 ), 
	.CO(\add_x_22_4/n1 ), 
	.B(\add_x_22_4/n2 ), 
	.A(\addr_calc/iir_read_calc/count[30] ));
   NAND2X1TS \add_x_22_4/U13  (.Y(\add_x_22_4/n10 ), 
	.B(\addr_calc/iir_read_calc/count[27] ), 
	.A(n1572));
   NAND2X1TS \add_x_22_4/U22  (.Y(\add_x_22_4/n17 ), 
	.B(n1926), 
	.A(\addr_calc/iir_read_calc/count[24] ));
   NAND2X1TS \add_x_22_4/U33  (.Y(\add_x_22_4/n26 ), 
	.B(\add_x_22_4/n27 ), 
	.A(\add_x_22_4/n43 ));
   NAND2X1TS \add_x_22_4/U35  (.Y(\add_x_22_4/n28 ), 
	.B(n2565), 
	.A(n2031));
   XNOR2X1TS \add_x_22_4/U62  (.Y(\addr_calc/iir_read_calc/counter/N60 ), 
	.B(n1919), 
	.A(\add_x_22_4/n54 ));
   NAND2X1TS \add_x_22_4/U44  (.Y(\add_x_22_4/n35 ), 
	.B(n1687), 
	.A(n2028));
   NAND2X1TS \add_x_22_4/U53  (.Y(\add_x_22_4/n42 ), 
	.B(\add_x_22_4/n43 ), 
	.A(FE_OFN150_add_x_22_4_n59));
   NAND2X1TS \add_x_22_4/U55  (.Y(\add_x_22_4/n44 ), 
	.B(\addr_calc/iir_read_calc/count[19] ), 
	.A(n2025));
   NAND2X1TS \add_x_22_4/U64  (.Y(\add_x_22_4/n51 ), 
	.B(n1920), 
	.A(\addr_calc/iir_read_calc/count[16] ));
   NAND2X1TS \add_x_22_4/U148  (.Y(\add_x_22_4/n119 ), 
	.B(\addr_calc/iir_read_calc/count[0] ), 
	.A(n1898));
   NAND2X1TS \add_x_22_4/U139  (.Y(\add_x_22_4/n112 ), 
	.B(\addr_calc/iir_read_calc/count[3] ), 
	.A(n2015));
   NAND2X1TS \add_x_22_4/U128  (.Y(\add_x_22_4/n103 ), 
	.B(\addr_calc/iir_read_calc/count[5] ), 
	.A(FE_OFN244_addr_calc_iir_read_calc_count_4_));
   NAND2X1TS \add_x_22_4/U86  (.Y(\add_x_22_4/n69 ), 
	.B(\addr_calc/iir_read_calc/count[13] ), 
	.A(\addr_calc/iir_read_calc/count[12] ));
   NAND2X1TS \add_x_22_4/U97  (.Y(\add_x_22_4/n78 ), 
	.B(FE_OFN236_addr_calc_iir_read_calc_count_11_), 
	.A(\addr_calc/iir_read_calc/count[10] ));
   NAND2X1TS \add_x_22_4/U108  (.Y(\add_x_22_4/n87 ), 
	.B(n1685), 
	.A(\addr_calc/iir_read_calc/count[8] ));
   XOR2X1TS \add_x_22_4/U136  (.Y(\addr_calc/iir_read_calc/counter/N46 ), 
	.B(n1901), 
	.A(\add_x_22_4/n115 ));
   XOR2X1TS \add_x_22_4/U115  (.Y(\addr_calc/iir_read_calc/counter/N50 ), 
	.B(\add_x_22_4/n98 ), 
	.A(\add_x_22_4/n99 ));
   XOR2X1TS \add_x_22_4/U105  (.Y(\addr_calc/iir_read_calc/counter/N52 ), 
	.B(n1907), 
	.A(\add_x_22_4/n90 ));
   XOR2X1TS \add_x_22_4/U100  (.Y(\addr_calc/iir_read_calc/counter/N53 ), 
	.B(\add_x_22_4/n84 ), 
	.A(\add_x_22_4/n85 ));
   XOR2X1TS \add_x_22_4/U72  (.Y(\addr_calc/iir_read_calc/counter/N58 ), 
	.B(\add_x_22_4/n64 ), 
	.A(\add_x_22_4/n65 ));
   XOR2X1TS \add_x_22_4/U67  (.Y(\addr_calc/iir_read_calc/counter/N59 ), 
	.B(\add_x_22_4/n57 ), 
	.A(\add_x_22_4/n58 ));
   XOR2X1TS \add_x_22_4/U51  (.Y(\addr_calc/iir_read_calc/counter/N62 ), 
	.B(\add_x_22_4/n46 ), 
	.A(\add_x_22_4/n47 ));
   XOR2X1TS \add_x_22_4/U20  (.Y(\addr_calc/iir_read_calc/counter/N68 ), 
	.B(n1925), 
	.A(\add_x_22_4/n20 ));
   XOR2X1TS \add_x_22_4/U4  (.Y(\addr_calc/iir_read_calc/counter/N71 ), 
	.B(\add_x_22_4/n7 ), 
	.A(\add_x_22_4/n8 ));
   XOR2X1TS \add_x_22_4/U1  (.Y(\addr_calc/iir_read_calc/counter/N74 ), 
	.B(\addr_calc/iir_read_calc/count[31] ), 
	.A(\add_x_22_4/n1 ));
   NOR2X1TS \add_x_22_1/U127  (.Y(\add_x_22_1/n102 ), 
	.B(\add_x_22_1/n103 ), 
	.A(\add_x_22_1/n110 ));
   NOR2X1TS \add_x_22_1/U85  (.Y(\add_x_22_1/n68 ), 
	.B(\add_x_22_1/n69 ), 
	.A(\add_x_22_1/n76 ));
   NOR2X1TS \add_x_22_1/U63  (.Y(\add_x_22_1/n50 ), 
	.B(\add_x_22_1/n51 ), 
	.A(\add_x_22_1/n58 ));
   NOR2X1TS \add_x_22_1/U68  (.Y(\add_x_22_1/n54 ), 
	.B(\add_x_22_1/n57 ), 
	.A(\add_x_22_1/n58 ));
   NOR2X1TS \add_x_22_1/U43  (.Y(\add_x_22_1/n34 ), 
	.B(\add_x_22_1/n35 ), 
	.A(\add_x_22_1/n42 ));
   NOR2X1TS \add_x_22_1/U21  (.Y(\add_x_22_1/n16 ), 
	.B(\add_x_22_1/n17 ), 
	.A(\add_x_22_1/n24 ));
   NOR2X1TS \add_x_22_1/U6  (.Y(\add_x_22_1/n4 ), 
	.B(\add_x_22_1/n5 ), 
	.A(\add_x_22_1/n26 ));
   NOR2X1TS \add_x_22_1/U12  (.Y(\add_x_22_1/n9 ), 
	.B(\add_x_22_1/n10 ), 
	.A(\add_x_22_1/n17 ));
   NOR2X1TS \add_x_22_1/U34  (.Y(\add_x_22_1/n27 ), 
	.B(\add_x_22_1/n28 ), 
	.A(\add_x_22_1/n35 ));
   NOR2X1TS \add_x_22_1/U54  (.Y(\add_x_22_1/n43 ), 
	.B(\add_x_22_1/n44 ), 
	.A(\add_x_22_1/n51 ));
   NOR2X1TS \add_x_22_1/U138  (.Y(\add_x_22_1/n111 ), 
	.B(\add_x_22_1/n119 ), 
	.A(\add_x_22_1/n112 ));
   NOR2X1TS \add_x_22_1/U118  (.Y(\add_x_22_1/n95 ), 
	.B(\add_x_22_1/n96 ), 
	.A(\add_x_22_1/n103 ));
   NOR2X1TS \add_x_22_1/U96  (.Y(\add_x_22_1/n77 ), 
	.B(\add_x_22_1/n78 ), 
	.A(\add_x_22_1/n87 ));
   NAND2X1TS \add_x_22_1/U90  (.Y(\add_x_22_1/n72 ), 
	.B(n2023), 
	.A(\add_x_22_1/n75 ));
   XNOR2X1TS \add_x_22_1/U89  (.Y(\addr_calc/fft_write_calc/counter/N55 ), 
	.B(\add_x_22_1/n74 ), 
	.A(\add_x_22_1/n75 ));
   NAND2X1TS \add_x_22_1/U123  (.Y(\add_x_22_1/n99 ), 
	.B(FE_OFN272_addr_calc_fft_write_calc_count_6_), 
	.A(\add_x_22_1/n102 ));
   XNOR2X1TS \add_x_22_1/U111  (.Y(\addr_calc/fft_write_calc/counter/N51 ), 
	.B(\add_x_22_1/n92 ), 
	.A(\add_x_22_1/n93 ));
   XNOR2X1TS \add_x_22_1/U80  (.Y(\addr_calc/fft_write_calc/counter/N57 ), 
	.B(\add_x_22_1/n67 ), 
	.A(\add_x_22_1/n68 ));
   NAND2X1TS \add_x_22_1/U143  (.Y(\add_x_22_1/n115 ), 
	.B(n2032), 
	.A(\add_x_22_1/n118 ));
   NAND2X1TS \add_x_22_1/U95  (.Y(\add_x_22_1/n76 ), 
	.B(\add_x_22_1/n77 ), 
	.A(\add_x_22_1/n93 ));
   NAND2X1TS \add_x_22_1/U48  (.Y(\add_x_22_1/n38 ), 
	.B(\addr_calc/fft_write_calc/count[20] ), 
	.A(\add_x_22_1/n41 ));
   XNOR2X1TS \add_x_22_1/U62  (.Y(\addr_calc/fft_write_calc/counter/N60 ), 
	.B(\add_x_22_1/n53 ), 
	.A(\add_x_22_1/n54 ));
   NAND2X1TS \add_x_22_1/U53  (.Y(\add_x_22_1/n42 ), 
	.B(\add_x_22_1/n43 ), 
	.A(\add_x_22_1/n59 ));
   NAND2X1TS \add_x_22_1/U26  (.Y(\add_x_22_1/n20 ), 
	.B(FE_OFN276_addr_calc_fft_write_calc_count_24_), 
	.A(\add_x_22_1/n23 ));
   NAND2X1TS \add_x_22_1/U11  (.Y(\add_x_22_1/n8 ), 
	.B(\add_x_22_1/n9 ), 
	.A(\add_x_22_1/n23 ));
   ADDHXLTS \add_x_22_1/U2  (.S(\addr_calc/fft_write_calc/counter/N73 ), 
	.CO(\add_x_22_1/n1 ), 
	.B(\add_x_22_1/n2 ), 
	.A(\addr_calc/fft_write_calc/count[30] ));
   NAND2X1TS \add_x_22_1/U22  (.Y(\add_x_22_1/n17 ), 
	.B(\addr_calc/fft_write_calc/count[25] ), 
	.A(FE_OFN277_addr_calc_fft_write_calc_count_24_));
   NAND2X1TS \add_x_22_1/U33  (.Y(\add_x_22_1/n26 ), 
	.B(\add_x_22_1/n27 ), 
	.A(\add_x_22_1/n43 ));
   NAND2X1TS \add_x_22_1/U35  (.Y(\add_x_22_1/n28 ), 
	.B(n2555), 
	.A(FE_OFN285_addr_calc_fft_write_calc_count_22_));
   NAND2X1TS \add_x_22_1/U44  (.Y(\add_x_22_1/n35 ), 
	.B(\addr_calc/fft_write_calc/count[21] ), 
	.A(\addr_calc/fft_write_calc/count[20] ));
   NAND2X1TS \add_x_22_1/U55  (.Y(\add_x_22_1/n44 ), 
	.B(\addr_calc/fft_write_calc/count[19] ), 
	.A(n2020));
   NAND2X1TS \add_x_22_1/U64  (.Y(\add_x_22_1/n51 ), 
	.B(n1924), 
	.A(n2567));
   NAND2X2TS \add_x_22_1/U117  (.Y(\add_x_22_1/n94 ), 
	.B(\add_x_22_1/n111 ), 
	.A(\add_x_22_1/n95 ));
   NAND2X1TS \add_x_22_1/U148  (.Y(\add_x_22_1/n119 ), 
	.B(FE_OFN260_addr_calc_fft_write_calc_count_0_), 
	.A(\addr_calc/fft_write_calc/count[1] ));
   NAND2X1TS \add_x_22_1/U139  (.Y(\add_x_22_1/n112 ), 
	.B(\addr_calc/fft_write_calc/count[3] ), 
	.A(\addr_calc/fft_write_calc/count[2] ));
   NAND2X1TS \add_x_22_1/U119  (.Y(\add_x_22_1/n96 ), 
	.B(\addr_calc/fft_write_calc/count[7] ), 
	.A(FE_OFN272_addr_calc_fft_write_calc_count_6_));
   NAND2X1TS \add_x_22_1/U86  (.Y(\add_x_22_1/n69 ), 
	.B(\addr_calc/fft_write_calc/count[13] ), 
	.A(\addr_calc/fft_write_calc/count[12] ));
   NAND2X1TS \add_x_22_1/U97  (.Y(\add_x_22_1/n78 ), 
	.B(\addr_calc/fft_write_calc/count[11] ), 
	.A(\addr_calc/fft_write_calc/count[10] ));
   NAND2X1TS \add_x_22_1/U108  (.Y(\add_x_22_1/n87 ), 
	.B(\addr_calc/fft_write_calc/count[9] ), 
	.A(\addr_calc/fft_write_calc/count[8] ));
   XOR2X1TS \add_x_22_1/U136  (.Y(\addr_calc/fft_write_calc/counter/N46 ), 
	.B(\add_x_22_1/n114 ), 
	.A(\add_x_22_1/n115 ));
   XOR2X1TS \add_x_22_1/U131  (.Y(\addr_calc/fft_write_calc/counter/N47 ), 
	.B(\add_x_22_1/n109 ), 
	.A(\add_x_22_1/n110 ));
   XOR2X1TS \add_x_22_1/U115  (.Y(\addr_calc/fft_write_calc/counter/N50 ), 
	.B(\add_x_22_1/n98 ), 
	.A(\add_x_22_1/n99 ));
   XOR2X1TS \add_x_22_1/U105  (.Y(\addr_calc/fft_write_calc/counter/N52 ), 
	.B(\add_x_22_1/n89 ), 
	.A(\add_x_22_1/n90 ));
   XOR2X1TS \add_x_22_1/U100  (.Y(\addr_calc/fft_write_calc/counter/N53 ), 
	.B(\add_x_22_1/n84 ), 
	.A(\add_x_22_1/n85 ));
   XOR2X1TS \add_x_22_1/U84  (.Y(\addr_calc/fft_write_calc/counter/N56 ), 
	.B(\add_x_22_1/n71 ), 
	.A(\add_x_22_1/n72 ));
   XOR2X1TS \add_x_22_1/U72  (.Y(\addr_calc/fft_write_calc/counter/N58 ), 
	.B(\add_x_22_1/n64 ), 
	.A(\add_x_22_1/n65 ));
   XOR2X1TS \add_x_22_1/U67  (.Y(\addr_calc/fft_write_calc/counter/N59 ), 
	.B(\add_x_22_1/n57 ), 
	.A(\add_x_22_1/n58 ));
   XOR2X1TS \add_x_22_1/U51  (.Y(\addr_calc/fft_write_calc/counter/N62 ), 
	.B(n1921), 
	.A(\add_x_22_1/n47 ));
   XOR2X1TS \add_x_22_1/U42  (.Y(\addr_calc/fft_write_calc/counter/N64 ), 
	.B(n1917), 
	.A(\add_x_22_1/n38 ));
   XOR2X1TS \add_x_22_1/U29  (.Y(\addr_calc/fft_write_calc/counter/N66 ), 
	.B(\add_x_22_1/n30 ), 
	.A(\add_x_22_1/n31 ));
   XOR2X1TS \add_x_22_1/U20  (.Y(\addr_calc/fft_write_calc/counter/N68 ), 
	.B(n1914), 
	.A(\add_x_22_1/n20 ));
   XOR2X1TS \add_x_22_1/U4  (.Y(\addr_calc/fft_write_calc/counter/N71 ), 
	.B(\add_x_22_1/n7 ), 
	.A(\add_x_22_1/n8 ));
   AHHCINX2TS \add_x_22_1/U3  (.S(\addr_calc/fft_write_calc/counter/N72 ), 
	.CO(\add_x_22_1/n2 ), 
	.CIN(\add_x_22_1/n3 ), 
	.A(\addr_calc/fft_write_calc/count[29] ));
   XOR2X1TS \add_x_22_1/U1  (.Y(\addr_calc/fft_write_calc/counter/N74 ), 
	.B(\addr_calc/fft_write_calc/count[31] ), 
	.A(\add_x_22_1/n1 ));
   NOR2X1TS \add_x_22_5/U101  (.Y(\add_x_22_5/n81 ), 
	.B(\add_x_22_5/n84 ), 
	.A(\add_x_22_5/n85 ));
   NOR2X1TS \add_x_22_5/U132  (.Y(\add_x_22_5/n106 ), 
	.B(\add_x_22_5/n109 ), 
	.A(\add_x_22_5/n110 ));
   NOR2X1TS \add_x_22_5/U127  (.Y(\add_x_22_5/n102 ), 
	.B(\add_x_22_5/n103 ), 
	.A(\add_x_22_5/n110 ));
   NOR2X1TS \add_x_22_5/U21  (.Y(\add_x_22_5/n16 ), 
	.B(\add_x_22_5/n17 ), 
	.A(\add_x_22_5/n24 ));
   NOR2X1TS \add_x_22_5/U85  (.Y(\add_x_22_5/n68 ), 
	.B(\add_x_22_5/n69 ), 
	.A(\add_x_22_5/n76 ));
   NOR2X1TS \add_x_22_5/U63  (.Y(\add_x_22_5/n50 ), 
	.B(\add_x_22_5/n51 ), 
	.A(\add_x_22_5/n58 ));
   NOR2X1TS \add_x_22_5/U43  (.Y(\add_x_22_5/n34 ), 
	.B(\add_x_22_5/n35 ), 
	.A(\add_x_22_5/n42 ));
   NOR2X1TS \add_x_22_5/U6  (.Y(\add_x_22_5/n4 ), 
	.B(\add_x_22_5/n5 ), 
	.A(\add_x_22_5/n26 ));
   NOR2X1TS \add_x_22_5/U12  (.Y(\add_x_22_5/n9 ), 
	.B(\add_x_22_5/n10 ), 
	.A(\add_x_22_5/n17 ));
   NOR2X1TS \add_x_22_5/U54  (.Y(\add_x_22_5/n43 ), 
	.B(\add_x_22_5/n44 ), 
	.A(\add_x_22_5/n51 ));
   NOR2X1TS \add_x_22_5/U68  (.Y(\add_x_22_5/n54 ), 
	.B(\add_x_22_5/n57 ), 
	.A(\add_x_22_5/n58 ));
   NOR2X1TS \add_x_22_5/U138  (.Y(\add_x_22_5/n111 ), 
	.B(\add_x_22_5/n119 ), 
	.A(\add_x_22_5/n112 ));
   NOR2X1TS \add_x_22_5/U96  (.Y(\add_x_22_5/n77 ), 
	.B(\add_x_22_5/n78 ), 
	.A(\add_x_22_5/n87 ));
   XNOR2X1TS \add_x_22_5/U146  (.Y(\addr_calc/iir_write_calc/counter/N44 ), 
	.B(n2578), 
	.A(\add_x_22_5/n121 ));
   XNOR2X1TS \add_x_22_5/U80  (.Y(\addr_calc/iir_write_calc/counter/N57 ), 
	.B(\add_x_22_5/n67 ), 
	.A(\add_x_22_5/n68 ));
   NAND2X1TS \add_x_22_5/U123  (.Y(\add_x_22_5/n99 ), 
	.B(n2039), 
	.A(\add_x_22_5/n102 ));
   XNOR2X1TS \add_x_22_5/U93  (.Y(\addr_calc/iir_write_calc/counter/N54 ), 
	.B(\add_x_22_5/n80 ), 
	.A(\add_x_22_5/n81 ));
   XNOR2X1TS \add_x_22_5/U126  (.Y(\addr_calc/iir_write_calc/counter/N48 ), 
	.B(n1937), 
	.A(\add_x_22_5/n106 ));
   XNOR2X1TS \add_x_22_5/U142  (.Y(\addr_calc/iir_write_calc/counter/N45 ), 
	.B(\add_x_22_5/n117 ), 
	.A(\add_x_22_5/n118 ));
   NAND2X1TS \add_x_22_5/U90  (.Y(\add_x_22_5/n72 ), 
	.B(n2044), 
	.A(\add_x_22_5/n75 ));
   XNOR2X1TS \add_x_22_5/U122  (.Y(\addr_calc/iir_write_calc/counter/N49 ), 
	.B(\add_x_22_5/n101 ), 
	.A(\add_x_22_5/n102 ));
   XNOR2X1TS \add_x_22_5/U111  (.Y(\addr_calc/iir_write_calc/counter/N51 ), 
	.B(\add_x_22_5/n92 ), 
	.A(\add_x_22_5/n93 ));
   XNOR2X1TS \add_x_22_5/U89  (.Y(\addr_calc/iir_write_calc/counter/N55 ), 
	.B(\add_x_22_5/n74 ), 
	.A(\add_x_22_5/n75 ));
   XNOR2X1TS \add_x_22_5/U16  (.Y(\addr_calc/iir_write_calc/counter/N69 ), 
	.B(\add_x_22_5/n15 ), 
	.A(\add_x_22_5/n16 ));
   NAND2X1TS \add_x_22_5/U17  (.Y(\add_x_22_5/n13 ), 
	.B(n2573), 
	.A(\add_x_22_5/n16 ));
   NAND2X1TS \add_x_22_5/U26  (.Y(\add_x_22_5/n20 ), 
	.B(\addr_calc/iir_write_calc/count[24] ), 
	.A(\add_x_22_5/n23 ));
   XNOR2X1TS \add_x_22_5/U25  (.Y(\addr_calc/iir_write_calc/counter/N67 ), 
	.B(n2050), 
	.A(\add_x_22_5/n23 ));
   NAND2X1TS \add_x_22_5/U11  (.Y(\add_x_22_5/n8 ), 
	.B(\add_x_22_5/n9 ), 
	.A(\add_x_22_5/n23 ));
   NAND2X1TS \add_x_22_5/U39  (.Y(\add_x_22_5/n31 ), 
	.B(n2579), 
	.A(\add_x_22_5/n34 ));
   NAND2X1TS \add_x_22_5/U95  (.Y(\add_x_22_5/n76 ), 
	.B(\add_x_22_5/n77 ), 
	.A(\add_x_22_5/n93 ));
   NAND2X1TS \add_x_22_5/U59  (.Y(\add_x_22_5/n47 ), 
	.B(FE_OFN266_addr_calc_iir_write_calc_count_18_), 
	.A(\add_x_22_5/n50 ));
   XNOR2X1TS \add_x_22_5/U38  (.Y(\addr_calc/iir_write_calc/counter/N65 ), 
	.B(\add_x_22_5/n33 ), 
	.A(\add_x_22_5/n34 ));
   NAND2X1TS \add_x_22_5/U53  (.Y(\add_x_22_5/n42 ), 
	.B(\add_x_22_5/n43 ), 
	.A(FE_OFN148_add_x_22_5_n59));
   ADDHXLTS \add_x_22_5/U2  (.S(\addr_calc/iir_write_calc/counter/N73 ), 
	.CO(\add_x_22_5/n1 ), 
	.B(\add_x_22_5/n2 ), 
	.A(FE_OFN239_addr_calc_iir_write_calc_count_30_));
   NAND2X1TS \add_x_22_5/U5  (.Y(\add_x_22_5/n3 ), 
	.B(FE_OFN148_add_x_22_5_n59), 
	.A(\add_x_22_5/n4 ));
   NAND2X1TS \add_x_22_5/U22  (.Y(\add_x_22_5/n17 ), 
	.B(n1969), 
	.A(n2051));
   NAND2X1TS \add_x_22_5/U44  (.Y(\add_x_22_5/n35 ), 
	.B(n1962), 
	.A(n2048));
   NAND2X1TS \add_x_22_5/U55  (.Y(\add_x_22_5/n44 ), 
	.B(n1958), 
	.A(FE_OFN266_addr_calc_iir_write_calc_count_18_));
   NAND2X1TS \add_x_22_5/U64  (.Y(\add_x_22_5/n51 ), 
	.B(\addr_calc/iir_write_calc/count[17] ), 
	.A(\addr_calc/iir_write_calc/count[16] ));
   XNOR2X1TS \add_x_22_5/U62  (.Y(\addr_calc/iir_write_calc/counter/N60 ), 
	.B(\add_x_22_5/n53 ), 
	.A(\add_x_22_5/n54 ));
   NAND2X1TS \add_x_22_5/U148  (.Y(\add_x_22_5/n119 ), 
	.B(\addr_calc/iir_write_calc/count[0] ), 
	.A(n1931));
   NAND2X1TS \add_x_22_5/U139  (.Y(\add_x_22_5/n112 ), 
	.B(\addr_calc/iir_write_calc/count[3] ), 
	.A(n2036));
   NAND2X1TS \add_x_22_5/U128  (.Y(\add_x_22_5/n103 ), 
	.B(\addr_calc/iir_write_calc/count[5] ), 
	.A(\addr_calc/iir_write_calc/count[4] ));
   NAND2X1TS \add_x_22_5/U86  (.Y(\add_x_22_5/n69 ), 
	.B(\addr_calc/iir_write_calc/count[13] ), 
	.A(\addr_calc/iir_write_calc/count[12] ));
   NAND2X1TS \add_x_22_5/U97  (.Y(\add_x_22_5/n78 ), 
	.B(\addr_calc/iir_write_calc/count[11] ), 
	.A(\addr_calc/iir_write_calc/count[10] ));
   NAND2X1TS \add_x_22_5/U108  (.Y(\add_x_22_5/n87 ), 
	.B(\addr_calc/iir_write_calc/count[9] ), 
	.A(\addr_calc/iir_write_calc/count[8] ));
   XOR2X1TS \add_x_22_5/U136  (.Y(\addr_calc/iir_write_calc/counter/N46 ), 
	.B(\add_x_22_5/n114 ), 
	.A(\add_x_22_5/n115 ));
   XOR2X1TS \add_x_22_5/U131  (.Y(\addr_calc/iir_write_calc/counter/N47 ), 
	.B(\add_x_22_5/n109 ), 
	.A(\add_x_22_5/n110 ));
   XOR2X1TS \add_x_22_5/U115  (.Y(\addr_calc/iir_write_calc/counter/N50 ), 
	.B(n1938), 
	.A(\add_x_22_5/n99 ));
   XOR2X1TS \add_x_22_5/U105  (.Y(\addr_calc/iir_write_calc/counter/N52 ), 
	.B(\add_x_22_5/n89 ), 
	.A(\add_x_22_5/n90 ));
   XOR2X1TS \add_x_22_5/U100  (.Y(\addr_calc/iir_write_calc/counter/N53 ), 
	.B(\add_x_22_5/n84 ), 
	.A(\add_x_22_5/n85 ));
   XOR2X1TS \add_x_22_5/U84  (.Y(\addr_calc/iir_write_calc/counter/N56 ), 
	.B(\add_x_22_5/n71 ), 
	.A(\add_x_22_5/n72 ));
   XOR2X1TS \add_x_22_5/U51  (.Y(\addr_calc/iir_write_calc/counter/N62 ), 
	.B(n1957), 
	.A(\add_x_22_5/n47 ));
   XOR2X1TS \add_x_22_5/U29  (.Y(\addr_calc/iir_write_calc/counter/N66 ), 
	.B(n1964), 
	.A(\add_x_22_5/n31 ));
   XOR2X1TS \add_x_22_5/U20  (.Y(\addr_calc/iir_write_calc/counter/N68 ), 
	.B(n1968), 
	.A(\add_x_22_5/n20 ));
   XOR2X1TS \add_x_22_5/U10  (.Y(\addr_calc/iir_write_calc/counter/N70 ), 
	.B(n1971), 
	.A(\add_x_22_5/n13 ));
   XOR2X1TS \add_x_22_5/U4  (.Y(\addr_calc/iir_write_calc/counter/N71 ), 
	.B(n1973), 
	.A(\add_x_22_5/n8 ));
   AHHCINX2TS \add_x_22_5/U3  (.S(\addr_calc/iir_write_calc/counter/N72 ), 
	.CO(\add_x_22_5/n2 ), 
	.CIN(\add_x_22_5/n3 ), 
	.A(n1851));
   XOR2X1TS \add_x_22_5/U1  (.Y(\addr_calc/iir_write_calc/counter/N74 ), 
	.B(FE_OFN240_addr_calc_iir_write_calc_count_31_), 
	.A(\add_x_22_5/n1 ));
   NOR2X1TS \add_x_22_3/U101  (.Y(\add_x_22_3/n81 ), 
	.B(\add_x_22_3/n84 ), 
	.A(\add_x_22_3/n85 ));
   NOR2X1TS \add_x_22_3/U132  (.Y(\add_x_22_3/n106 ), 
	.B(\add_x_22_3/n109 ), 
	.A(\add_x_22_3/n110 ));
   NOR2X1TS \add_x_22_3/U127  (.Y(\add_x_22_3/n102 ), 
	.B(\add_x_22_3/n103 ), 
	.A(\add_x_22_3/n110 ));
   NOR2X1TS \add_x_22_3/U63  (.Y(\add_x_22_3/n50 ), 
	.B(\add_x_22_3/n51 ), 
	.A(\add_x_22_3/n58 ));
   NOR2X1TS \add_x_22_3/U85  (.Y(\add_x_22_3/n68 ), 
	.B(\add_x_22_3/n69 ), 
	.A(\add_x_22_3/n76 ));
   NOR2X1TS \add_x_22_3/U43  (.Y(\add_x_22_3/n34 ), 
	.B(\add_x_22_3/n35 ), 
	.A(\add_x_22_3/n42 ));
   NOR2X1TS \add_x_22_3/U21  (.Y(\add_x_22_3/n16 ), 
	.B(\add_x_22_3/n17 ), 
	.A(\add_x_22_3/n24 ));
   NOR2X1TS \add_x_22_3/U12  (.Y(\add_x_22_3/n9 ), 
	.B(\add_x_22_3/n10 ), 
	.A(\add_x_22_3/n17 ));
   NOR2X1TS \add_x_22_3/U34  (.Y(\add_x_22_3/n27 ), 
	.B(\add_x_22_3/n28 ), 
	.A(\add_x_22_3/n35 ));
   NOR2X1TS \add_x_22_3/U54  (.Y(\add_x_22_3/n43 ), 
	.B(\add_x_22_3/n44 ), 
	.A(\add_x_22_3/n51 ));
   NOR2X1TS \add_x_22_3/U68  (.Y(\add_x_22_3/n54 ), 
	.B(\add_x_22_3/n57 ), 
	.A(\add_x_22_3/n58 ));
   NOR2X1TS \add_x_22_3/U138  (.Y(\add_x_22_3/n111 ), 
	.B(\add_x_22_3/n119 ), 
	.A(\add_x_22_3/n112 ));
   NOR2X1TS \add_x_22_3/U96  (.Y(\add_x_22_3/n77 ), 
	.B(\add_x_22_3/n78 ), 
	.A(\add_x_22_3/n87 ));
   XNOR2X1TS \add_x_22_3/U142  (.Y(\addr_calc/fir_write_calc/counter/N45 ), 
	.B(n1989), 
	.A(\add_x_22_3/n118 ));
   NAND2X1TS \add_x_22_3/U143  (.Y(\add_x_22_3/n115 ), 
	.B(\addr_calc/fir_write_calc/count[2] ), 
	.A(\add_x_22_3/n118 ));
   XNOR2X1TS \add_x_22_3/U111  (.Y(\addr_calc/fir_write_calc/counter/N51 ), 
	.B(\add_x_22_3/n92 ), 
	.A(\add_x_22_3/n93 ));
   XNOR2X1TS \add_x_22_3/U93  (.Y(\addr_calc/fir_write_calc/counter/N54 ), 
	.B(\add_x_22_3/n80 ), 
	.A(\add_x_22_3/n81 ));
   XNOR2X1TS \add_x_22_3/U126  (.Y(\addr_calc/fir_write_calc/counter/N48 ), 
	.B(\add_x_22_3/n105 ), 
	.A(\add_x_22_3/n106 ));
   XNOR2X1TS \add_x_22_3/U38  (.Y(\addr_calc/fir_write_calc/counter/N65 ), 
	.B(n2012), 
	.A(\add_x_22_3/n34 ));
   XNOR2X1TS \add_x_22_3/U122  (.Y(\addr_calc/fir_write_calc/counter/N49 ), 
	.B(\add_x_22_3/n101 ), 
	.A(\add_x_22_3/n102 ));
   XNOR2X1TS \add_x_22_3/U80  (.Y(\addr_calc/fir_write_calc/counter/N57 ), 
	.B(n2002), 
	.A(\add_x_22_3/n68 ));
   XNOR2X1TS \add_x_22_3/U58  (.Y(\addr_calc/fir_write_calc/counter/N61 ), 
	.B(n2005), 
	.A(\add_x_22_3/n50 ));
   NAND2X1TS \add_x_22_3/U90  (.Y(\add_x_22_3/n72 ), 
	.B(FE_OFN233_addr_calc_fir_write_calc_count_12_), 
	.A(\add_x_22_3/n75 ));
   NAND2X1TS \add_x_22_3/U59  (.Y(\add_x_22_3/n47 ), 
	.B(n2006), 
	.A(\add_x_22_3/n50 ));
   NAND2X1TS \add_x_22_3/U95  (.Y(\add_x_22_3/n76 ), 
	.B(\add_x_22_3/n77 ), 
	.A(\add_x_22_3/n93 ));
   NAND2X1TS \add_x_22_3/U17  (.Y(\add_x_22_3/n13 ), 
	.B(FE_OFN268_addr_calc_fir_write_calc_count_26_), 
	.A(\add_x_22_3/n16 ));
   NAND2X1TS \add_x_22_3/U39  (.Y(\add_x_22_3/n31 ), 
	.B(n1668), 
	.A(\add_x_22_3/n34 ));
   NAND2X1TS \add_x_22_3/U53  (.Y(\add_x_22_3/n42 ), 
	.B(\add_x_22_3/n43 ), 
	.A(\add_x_22_3/n59 ));
   NAND2X1TS \add_x_22_3/U11  (.Y(\add_x_22_3/n8 ), 
	.B(\add_x_22_3/n9 ), 
	.A(\add_x_22_3/n23 ));
   ADDHXLTS \add_x_22_3/U2  (.S(\addr_calc/fir_write_calc/counter/N73 ), 
	.CO(\add_x_22_3/n1 ), 
	.B(\add_x_22_3/n2 ), 
	.A(FE_OFN238_addr_calc_fir_write_calc_count_30_));
   NAND2X1TS \add_x_22_3/U22  (.Y(\add_x_22_3/n17 ), 
	.B(\addr_calc/fir_write_calc/count[25] ), 
	.A(n2577));
   NAND2X1TS \add_x_22_3/U26  (.Y(\add_x_22_3/n20 ), 
	.B(n2577), 
	.A(\add_x_22_3/n23 ));
   XNOR2X1TS \add_x_22_3/U25  (.Y(\addr_calc/fir_write_calc/counter/N67 ), 
	.B(\add_x_22_3/n22 ), 
	.A(\add_x_22_3/n23 ));
   NAND2X1TS \add_x_22_3/U33  (.Y(\add_x_22_3/n26 ), 
	.B(\add_x_22_3/n27 ), 
	.A(\add_x_22_3/n43 ));
   NAND2X1TS \add_x_22_3/U44  (.Y(\add_x_22_3/n35 ), 
	.B(n1892), 
	.A(FE_OFN282_addr_calc_fir_write_calc_count_20_));
   NAND2X1TS \add_x_22_3/U55  (.Y(\add_x_22_3/n44 ), 
	.B(n1670), 
	.A(n2006));
   NAND2X1TS \add_x_22_3/U64  (.Y(\add_x_22_3/n51 ), 
	.B(\addr_calc/fir_write_calc/count[17] ), 
	.A(n2564));
   XNOR2X1TS \add_x_22_3/U62  (.Y(\addr_calc/fir_write_calc/counter/N60 ), 
	.B(n1885), 
	.A(\add_x_22_3/n54 ));
   NAND2X1TS \add_x_22_3/U148  (.Y(\add_x_22_3/n119 ), 
	.B(FE_OFN252_addr_calc_fir_write_calc_count_0_), 
	.A(FE_OFN242_addr_calc_fir_write_calc_count_1_));
   NAND2X1TS \add_x_22_3/U139  (.Y(\add_x_22_3/n112 ), 
	.B(\addr_calc/fir_write_calc/count[3] ), 
	.A(n1990));
   NAND2X1TS \add_x_22_3/U128  (.Y(\add_x_22_3/n103 ), 
	.B(n1867), 
	.A(\addr_calc/fir_write_calc/count[4] ));
   NAND2X1TS \add_x_22_3/U86  (.Y(\add_x_22_3/n69 ), 
	.B(n1880), 
	.A(FE_OFN232_addr_calc_fir_write_calc_count_12_));
   NAND2X1TS \add_x_22_3/U97  (.Y(\add_x_22_3/n78 ), 
	.B(\addr_calc/fir_write_calc/count[11] ), 
	.A(n1874));
   NAND2X1TS \add_x_22_3/U108  (.Y(\add_x_22_3/n87 ), 
	.B(\addr_calc/fir_write_calc/count[9] ), 
	.A(FE_OFN257_addr_calc_fir_write_calc_count_8_));
   XOR2X1TS \add_x_22_3/U136  (.Y(\addr_calc/fir_write_calc/counter/N46 ), 
	.B(\add_x_22_3/n114 ), 
	.A(\add_x_22_3/n115 ));
   XOR2X1TS \add_x_22_3/U105  (.Y(\addr_calc/fir_write_calc/counter/N52 ), 
	.B(\add_x_22_3/n89 ), 
	.A(\add_x_22_3/n90 ));
   XOR2X1TS \add_x_22_3/U84  (.Y(\addr_calc/fir_write_calc/counter/N56 ), 
	.B(\add_x_22_3/n71 ), 
	.A(\add_x_22_3/n72 ));
   XOR2X1TS \add_x_22_3/U67  (.Y(\addr_calc/fir_write_calc/counter/N59 ), 
	.B(\add_x_22_3/n57 ), 
	.A(\add_x_22_3/n58 ));
   XOR2X1TS \add_x_22_3/U51  (.Y(\addr_calc/fir_write_calc/counter/N62 ), 
	.B(n1889), 
	.A(\add_x_22_3/n47 ));
   XOR2X1TS \add_x_22_3/U29  (.Y(\addr_calc/fir_write_calc/counter/N66 ), 
	.B(\add_x_22_3/n30 ), 
	.A(\add_x_22_3/n31 ));
   XOR2X1TS \add_x_22_3/U20  (.Y(\addr_calc/fir_write_calc/counter/N68 ), 
	.B(\add_x_22_3/n19 ), 
	.A(\add_x_22_3/n20 ));
   XOR2X1TS \add_x_22_3/U10  (.Y(\addr_calc/fir_write_calc/counter/N70 ), 
	.B(n1834), 
	.A(\add_x_22_3/n13 ));
   XOR2X1TS \add_x_22_3/U4  (.Y(\addr_calc/fir_write_calc/counter/N71 ), 
	.B(\add_x_22_3/n7 ), 
	.A(\add_x_22_3/n8 ));
   XOR2X1TS \add_x_22_3/U1  (.Y(\addr_calc/fir_write_calc/counter/N74 ), 
	.B(\addr_calc/fir_write_calc/count[31] ), 
	.A(\add_x_22_3/n1 ));
   NOR2X1TS \add_x_22_2/U68  (.Y(\add_x_22_2/n54 ), 
	.B(n1887), 
	.A(\add_x_22_2/n58 ));
   NOR2X1TS \add_x_22_2/U127  (.Y(\add_x_22_2/n102 ), 
	.B(\add_x_22_2/n103 ), 
	.A(\add_x_22_2/n110 ));
   NOR2X1TS \add_x_22_2/U101  (.Y(\add_x_22_2/n81 ), 
	.B(n1897), 
	.A(\add_x_22_2/n85 ));
   NOR2X1TS \add_x_22_2/U85  (.Y(\add_x_22_2/n68 ), 
	.B(\add_x_22_2/n69 ), 
	.A(\add_x_22_2/n76 ));
   NOR2X1TS \add_x_22_2/U63  (.Y(\add_x_22_2/n50 ), 
	.B(\add_x_22_2/n51 ), 
	.A(\add_x_22_2/n58 ));
   NOR2X1TS \add_x_22_2/U43  (.Y(\add_x_22_2/n34 ), 
	.B(\add_x_22_2/n35 ), 
	.A(\add_x_22_2/n42 ));
   NOR2X1TS \add_x_22_2/U12  (.Y(\add_x_22_2/n9 ), 
	.B(\add_x_22_2/n10 ), 
	.A(\add_x_22_2/n17 ));
   NOR2X1TS \add_x_22_2/U21  (.Y(\add_x_22_2/n16 ), 
	.B(\add_x_22_2/n17 ), 
	.A(\add_x_22_2/n24 ));
   NOR2X1TS \add_x_22_2/U54  (.Y(\add_x_22_2/n43 ), 
	.B(\add_x_22_2/n44 ), 
	.A(\add_x_22_2/n51 ));
   NOR2X1TS \add_x_22_2/U138  (.Y(\add_x_22_2/n111 ), 
	.B(\add_x_22_2/n119 ), 
	.A(\add_x_22_2/n112 ));
   NOR2X1TS \add_x_22_2/U96  (.Y(\add_x_22_2/n77 ), 
	.B(\add_x_22_2/n78 ), 
	.A(\add_x_22_2/n87 ));
   XNOR2X1TS \add_x_22_2/U142  (.Y(\addr_calc/fir_read_calc/counter/N45 ), 
	.B(\add_x_22_2/n117 ), 
	.A(\add_x_22_2/n118 ));
   XNOR2X1TS \add_x_22_2/U58  (.Y(\addr_calc/fir_read_calc/counter/N61 ), 
	.B(n1987), 
	.A(\add_x_22_2/n50 ));
   XNOR2X1TS \add_x_22_2/U89  (.Y(\addr_calc/fir_read_calc/counter/N55 ), 
	.B(\add_x_22_2/n74 ), 
	.A(\add_x_22_2/n75 ));
   XNOR2X1TS \add_x_22_2/U122  (.Y(\addr_calc/fir_read_calc/counter/N49 ), 
	.B(\add_x_22_2/n101 ), 
	.A(\add_x_22_2/n102 ));
   XNOR2X1TS \add_x_22_2/U62  (.Y(\addr_calc/fir_read_calc/counter/N60 ), 
	.B(\add_x_22_2/n53 ), 
	.A(\add_x_22_2/n54 ));
   XNOR2X1TS \add_x_22_2/U126  (.Y(\addr_calc/fir_read_calc/counter/N48 ), 
	.B(\add_x_22_2/n105 ), 
	.A(\add_x_22_2/n106 ));
   XNOR2X1TS \add_x_22_2/U47  (.Y(\addr_calc/fir_read_calc/counter/N63 ), 
	.B(n1984), 
	.A(\add_x_22_2/n41 ));
   NAND2X1TS \add_x_22_2/U90  (.Y(\add_x_22_2/n72 ), 
	.B(n1994), 
	.A(\add_x_22_2/n75 ));
   XNOR2X1TS \add_x_22_2/U80  (.Y(\addr_calc/fir_read_calc/counter/N57 ), 
	.B(n1991), 
	.A(\add_x_22_2/n68 ));
   NAND2X1TS \add_x_22_2/U48  (.Y(\add_x_22_2/n38 ), 
	.B(\addr_calc/fir_read_calc/count[20] ), 
	.A(\add_x_22_2/n41 ));
   XNOR2X1TS \add_x_22_2/U93  (.Y(\addr_calc/fir_read_calc/counter/N54 ), 
	.B(\add_x_22_2/n80 ), 
	.A(\add_x_22_2/n81 ));
   NAND2X1TS \add_x_22_2/U95  (.Y(\add_x_22_2/n76 ), 
	.B(\add_x_22_2/n77 ), 
	.A(\add_x_22_2/n93 ));
   XNOR2X1TS \add_x_22_2/U38  (.Y(\addr_calc/fir_read_calc/counter/N65 ), 
	.B(n1981), 
	.A(\add_x_22_2/n34 ));
   XNOR2X1TS \add_x_22_2/U111  (.Y(\addr_calc/fir_read_calc/counter/N51 ), 
	.B(\add_x_22_2/n92 ), 
	.A(\add_x_22_2/n93 ));
   NAND2X1TS \add_x_22_2/U59  (.Y(\add_x_22_2/n47 ), 
	.B(\addr_calc/fir_read_calc/count[18] ), 
	.A(\add_x_22_2/n50 ));
   XNOR2X1TS \add_x_22_2/U25  (.Y(\addr_calc/fir_read_calc/counter/N67 ), 
	.B(n1982), 
	.A(\add_x_22_2/n23 ));
   NAND2X1TS \add_x_22_2/U39  (.Y(\add_x_22_2/n31 ), 
	.B(n1691), 
	.A(\add_x_22_2/n34 ));
   NAND2X1TS \add_x_22_2/U53  (.Y(\add_x_22_2/n42 ), 
	.B(\add_x_22_2/n43 ), 
	.A(FE_OFN147_add_x_22_2_n59));
   ADDHXLTS \add_x_22_2/U2  (.S(\addr_calc/fir_read_calc/counter/N73 ), 
	.CO(\add_x_22_2/n1 ), 
	.B(\add_x_22_2/n2 ), 
	.A(\addr_calc/fir_read_calc/count[30] ));
   NAND2X1TS \add_x_22_2/U11  (.Y(\add_x_22_2/n8 ), 
	.B(\add_x_22_2/n9 ), 
	.A(\add_x_22_2/n23 ));
   NAND2X1TS \add_x_22_2/U22  (.Y(\add_x_22_2/n17 ), 
	.B(\addr_calc/fir_read_calc/count[25] ), 
	.A(\addr_calc/fir_read_calc/count[24] ));
   NAND2X1TS \add_x_22_2/U44  (.Y(\add_x_22_2/n35 ), 
	.B(n1879), 
	.A(\addr_calc/fir_read_calc/count[20] ));
   NAND2X1TS \add_x_22_2/U55  (.Y(\add_x_22_2/n44 ), 
	.B(n1881), 
	.A(\addr_calc/fir_read_calc/count[18] ));
   NAND2X1TS \add_x_22_2/U64  (.Y(\add_x_22_2/n51 ), 
	.B(n1884), 
	.A(n1888));
   NAND2X1TS \add_x_22_2/U148  (.Y(\add_x_22_2/n119 ), 
	.B(\addr_calc/fir_read_calc/count[0] ), 
	.A(FE_OFN249_addr_calc_fir_read_calc_count_1_));
   NAND2X1TS \add_x_22_2/U139  (.Y(\add_x_22_2/n112 ), 
	.B(\addr_calc/fir_read_calc/count[3] ), 
	.A(\addr_calc/fir_read_calc/count[2] ));
   NAND2X1TS \add_x_22_2/U128  (.Y(\add_x_22_2/n103 ), 
	.B(FE_OFN245_addr_calc_fir_read_calc_count_5_), 
	.A(n1906));
   NAND2X1TS \add_x_22_2/U86  (.Y(\add_x_22_2/n69 ), 
	.B(n1893), 
	.A(\addr_calc/fir_read_calc/count[12] ));
   NAND2X1TS \add_x_22_2/U97  (.Y(\add_x_22_2/n78 ), 
	.B(\addr_calc/fir_read_calc/count[11] ), 
	.A(n1540));
   NAND2X1TS \add_x_22_2/U108  (.Y(\add_x_22_2/n87 ), 
	.B(n1900), 
	.A(\addr_calc/fir_read_calc/count[8] ));
   XOR2X1TS \add_x_22_2/U131  (.Y(\addr_calc/fir_read_calc/counter/N47 ), 
	.B(\add_x_22_2/n109 ), 
	.A(\add_x_22_2/n110 ));
   XOR2X1TS \add_x_22_2/U115  (.Y(\addr_calc/fir_read_calc/counter/N50 ), 
	.B(\add_x_22_2/n98 ), 
	.A(\add_x_22_2/n99 ));
   XOR2X1TS \add_x_22_2/U105  (.Y(\addr_calc/fir_read_calc/counter/N52 ), 
	.B(n1899), 
	.A(\add_x_22_2/n90 ));
   XOR2X1TS \add_x_22_2/U100  (.Y(\addr_calc/fir_read_calc/counter/N53 ), 
	.B(n1897), 
	.A(\add_x_22_2/n85 ));
   XOR2X1TS \add_x_22_2/U84  (.Y(\addr_calc/fir_read_calc/counter/N56 ), 
	.B(\add_x_22_2/n71 ), 
	.A(\add_x_22_2/n72 ));
   XOR2X1TS \add_x_22_2/U67  (.Y(\addr_calc/fir_read_calc/counter/N59 ), 
	.B(n1887), 
	.A(\add_x_22_2/n58 ));
   XOR2X1TS \add_x_22_2/U51  (.Y(\addr_calc/fir_read_calc/counter/N62 ), 
	.B(\add_x_22_2/n46 ), 
	.A(\add_x_22_2/n47 ));
   XOR2X1TS \add_x_22_2/U42  (.Y(\addr_calc/fir_read_calc/counter/N64 ), 
	.B(n1878), 
	.A(\add_x_22_2/n38 ));
   XOR2X1TS \add_x_22_2/U29  (.Y(\addr_calc/fir_read_calc/counter/N66 ), 
	.B(\add_x_22_2/n30 ), 
	.A(\add_x_22_2/n31 ));
   XOR2X1TS \add_x_22_2/U4  (.Y(\addr_calc/fir_read_calc/counter/N71 ), 
	.B(n1870), 
	.A(\add_x_22_2/n8 ));
   NOR2X1TS \add_x_22_0/U127  (.Y(\add_x_22_0/n102 ), 
	.B(\add_x_22_0/n103 ), 
	.A(\add_x_22_0/n110 ));
   NOR2X1TS \add_x_22_0/U132  (.Y(\add_x_22_0/n106 ), 
	.B(\add_x_22_0/n109 ), 
	.A(\add_x_22_0/n110 ));
   NOR2X1TS \add_x_22_0/U85  (.Y(\add_x_22_0/n68 ), 
	.B(\add_x_22_0/n69 ), 
	.A(\add_x_22_0/n76 ));
   NOR2X1TS \add_x_22_0/U21  (.Y(\add_x_22_0/n16 ), 
	.B(\add_x_22_0/n17 ), 
	.A(\add_x_22_0/n24 ));
   NOR2X1TS \add_x_22_0/U43  (.Y(\add_x_22_0/n34 ), 
	.B(\add_x_22_0/n35 ), 
	.A(\add_x_22_0/n42 ));
   NOR2X1TS \add_x_22_0/U6  (.Y(\add_x_22_0/n4 ), 
	.B(\add_x_22_0/n5 ), 
	.A(\add_x_22_0/n26 ));
   NOR2X1TS \add_x_22_0/U12  (.Y(\add_x_22_0/n9 ), 
	.B(\add_x_22_0/n10 ), 
	.A(\add_x_22_0/n17 ));
   NOR2X1TS \add_x_22_0/U54  (.Y(\add_x_22_0/n43 ), 
	.B(\add_x_22_0/n44 ), 
	.A(\add_x_22_0/n51 ));
   NOR2X1TS \add_x_22_0/U63  (.Y(\add_x_22_0/n50 ), 
	.B(\add_x_22_0/n51 ), 
	.A(\add_x_22_0/n58 ));
   NOR2X1TS \add_x_22_0/U138  (.Y(\add_x_22_0/n111 ), 
	.B(\add_x_22_0/n119 ), 
	.A(\add_x_22_0/n112 ));
   NOR2X1TS \add_x_22_0/U118  (.Y(\add_x_22_0/n95 ), 
	.B(\add_x_22_0/n96 ), 
	.A(\add_x_22_0/n103 ));
   NOR2X1TS \add_x_22_0/U96  (.Y(\add_x_22_0/n77 ), 
	.B(\add_x_22_0/n78 ), 
	.A(\add_x_22_0/n87 ));
   XNOR2X1TS \add_x_22_0/U146  (.Y(\addr_calc/fft_read_calc/counter/N44 ), 
	.B(FE_OFN517_addr_calc_fft_read_calc_count_0_), 
	.A(\add_x_22_0/n121 ));
   XNOR2X1TS \add_x_22_0/U142  (.Y(\addr_calc/fft_read_calc/counter/N45 ), 
	.B(\add_x_22_0/n117 ), 
	.A(\add_x_22_0/n118 ));
   XNOR2X1TS \add_x_22_0/U89  (.Y(\addr_calc/fft_read_calc/counter/N55 ), 
	.B(n2045), 
	.A(\add_x_22_0/n75 ));
   XNOR2X1TS \add_x_22_0/U47  (.Y(\addr_calc/fft_read_calc/counter/N63 ), 
	.B(\add_x_22_0/n40 ), 
	.A(\add_x_22_0/n41 ));
   NAND2X1TS \add_x_22_0/U143  (.Y(\add_x_22_0/n115 ), 
	.B(n2056), 
	.A(\add_x_22_0/n118 ));
   XNOR2X1TS \add_x_22_0/U80  (.Y(\addr_calc/fft_read_calc/counter/N57 ), 
	.B(n2042), 
	.A(\add_x_22_0/n68 ));
   XNOR2X1TS \add_x_22_0/U38  (.Y(\addr_calc/fft_read_calc/counter/N65 ), 
	.B(n2040), 
	.A(\add_x_22_0/n34 ));
   XNOR2X1TS \add_x_22_0/U111  (.Y(\addr_calc/fft_read_calc/counter/N51 ), 
	.B(\add_x_22_0/n92 ), 
	.A(\add_x_22_0/n93 ));
   NAND2X1TS \add_x_22_0/U90  (.Y(\add_x_22_0/n72 ), 
	.B(\addr_calc/fft_read_calc/count[12] ), 
	.A(\add_x_22_0/n75 ));
   XNOR2X1TS \add_x_22_0/U126  (.Y(\addr_calc/fft_read_calc/counter/N48 ), 
	.B(\add_x_22_0/n105 ), 
	.A(\add_x_22_0/n106 ));
   NAND2X1TS \add_x_22_0/U95  (.Y(\add_x_22_0/n76 ), 
	.B(\add_x_22_0/n77 ), 
	.A(\add_x_22_0/n93 ));
   NAND2X1TS \add_x_22_0/U26  (.Y(\add_x_22_0/n20 ), 
	.B(\addr_calc/fft_read_calc/count[24] ), 
	.A(\add_x_22_0/n23 ));
   NAND2X1TS \add_x_22_0/U11  (.Y(\add_x_22_0/n8 ), 
	.B(\add_x_22_0/n9 ), 
	.A(\add_x_22_0/n23 ));
   NAND2X1TS \add_x_22_0/U17  (.Y(\add_x_22_0/n13 ), 
	.B(n2575), 
	.A(\add_x_22_0/n16 ));
   NAND2X1TS \add_x_22_0/U39  (.Y(\add_x_22_0/n31 ), 
	.B(n1665), 
	.A(\add_x_22_0/n34 ));
   NAND2X1TS \add_x_22_0/U53  (.Y(\add_x_22_0/n42 ), 
	.B(\add_x_22_0/n43 ), 
	.A(\add_x_22_0/n59 ));
   XNOR2X1TS \add_x_22_0/U25  (.Y(\addr_calc/fft_read_calc/counter/N67 ), 
	.B(n2037), 
	.A(\add_x_22_0/n23 ));
   ADDHXLTS \add_x_22_0/U2  (.S(\addr_calc/fft_read_calc/counter/N73 ), 
	.CO(\add_x_22_0/n1 ), 
	.B(\add_x_22_0/n2 ), 
	.A(\addr_calc/fft_read_calc/count[30] ));
   NAND2X1TS \add_x_22_0/U5  (.Y(\add_x_22_0/n3 ), 
	.B(\add_x_22_0/n59 ), 
	.A(\add_x_22_0/n4 ));
   NAND2X1TS \add_x_22_0/U7  (.Y(\add_x_22_0/n5 ), 
	.B(n2559), 
	.A(\add_x_22_0/n9 ));
   NAND2X1TS \add_x_22_0/U22  (.Y(\add_x_22_0/n17 ), 
	.B(\addr_calc/fft_read_calc/count[25] ), 
	.A(\addr_calc/fft_read_calc/count[24] ));
   NAND2X1TS \add_x_22_0/U44  (.Y(\add_x_22_0/n35 ), 
	.B(\addr_calc/fft_read_calc/count[21] ), 
	.A(n2572));
   NAND2X1TS \add_x_22_0/U55  (.Y(\add_x_22_0/n44 ), 
	.B(\addr_calc/fft_read_calc/count[19] ), 
	.A(n2569));
   NAND2X1TS \add_x_22_0/U59  (.Y(\add_x_22_0/n47 ), 
	.B(n2569), 
	.A(\add_x_22_0/n50 ));
   NAND2X1TS \add_x_22_0/U64  (.Y(\add_x_22_0/n51 ), 
	.B(\addr_calc/fft_read_calc/count[17] ), 
	.A(n2554));
   NAND2X2TS \add_x_22_0/U117  (.Y(\add_x_22_0/n94 ), 
	.B(\add_x_22_0/n111 ), 
	.A(\add_x_22_0/n95 ));
   NAND2X1TS \add_x_22_0/U148  (.Y(\add_x_22_0/n119 ), 
	.B(n2058), 
	.A(n1979));
   NAND2X1TS \add_x_22_0/U139  (.Y(\add_x_22_0/n112 ), 
	.B(\addr_calc/fft_read_calc/count[3] ), 
	.A(n2056));
   NAND2X1TS \add_x_22_0/U119  (.Y(\add_x_22_0/n96 ), 
	.B(\addr_calc/fft_read_calc/count[7] ), 
	.A(FE_OFN224_addr_calc_fft_read_calc_count_6_));
   NAND2X1TS \add_x_22_0/U128  (.Y(\add_x_22_0/n103 ), 
	.B(\addr_calc/fft_read_calc/count[5] ), 
	.A(FE_OFN263_addr_calc_fft_read_calc_count_4_));
   NAND2X1TS \add_x_22_0/U86  (.Y(\add_x_22_0/n69 ), 
	.B(n1967), 
	.A(n2046));
   NAND2X1TS \add_x_22_0/U97  (.Y(\add_x_22_0/n78 ), 
	.B(\addr_calc/fft_read_calc/count[11] ), 
	.A(\addr_calc/fft_read_calc/count[10] ));
   NAND2X1TS \add_x_22_0/U108  (.Y(\add_x_22_0/n87 ), 
	.B(\addr_calc/fft_read_calc/count[9] ), 
	.A(\addr_calc/fft_read_calc/count[8] ));
   XOR2X1TS \add_x_22_0/U136  (.Y(\addr_calc/fft_read_calc/counter/N46 ), 
	.B(\add_x_22_0/n114 ), 
	.A(\add_x_22_0/n115 ));
   XOR2X1TS \add_x_22_0/U115  (.Y(\addr_calc/fft_read_calc/counter/N50 ), 
	.B(n1975), 
	.A(\add_x_22_0/n99 ));
   XOR2X1TS \add_x_22_0/U105  (.Y(\addr_calc/fft_read_calc/counter/N52 ), 
	.B(\add_x_22_0/n89 ), 
	.A(\add_x_22_0/n90 ));
   XOR2X1TS \add_x_22_0/U100  (.Y(\addr_calc/fft_read_calc/counter/N53 ), 
	.B(\add_x_22_0/n84 ), 
	.A(\add_x_22_0/n85 ));
   XOR2X1TS \add_x_22_0/U84  (.Y(\addr_calc/fft_read_calc/counter/N56 ), 
	.B(n1966), 
	.A(\add_x_22_0/n72 ));
   XOR2X1TS \add_x_22_0/U72  (.Y(\addr_calc/fft_read_calc/counter/N58 ), 
	.B(n1963), 
	.A(\add_x_22_0/n65 ));
   XOR2X1TS \add_x_22_0/U51  (.Y(\addr_calc/fft_read_calc/counter/N62 ), 
	.B(n1955), 
	.A(\add_x_22_0/n47 ));
   XOR2X1TS \add_x_22_0/U29  (.Y(\addr_calc/fft_read_calc/counter/N66 ), 
	.B(n1949), 
	.A(\add_x_22_0/n31 ));
   XOR2X1TS \add_x_22_0/U20  (.Y(\addr_calc/fft_read_calc/counter/N68 ), 
	.B(n1946), 
	.A(\add_x_22_0/n20 ));
   XOR2X1TS \add_x_22_0/U10  (.Y(\addr_calc/fft_read_calc/counter/N70 ), 
	.B(n1943), 
	.A(\add_x_22_0/n13 ));
   XOR2X1TS \add_x_22_0/U4  (.Y(\addr_calc/fft_read_calc/counter/N71 ), 
	.B(\add_x_22_0/n7 ), 
	.A(\add_x_22_0/n8 ));
   AHHCINX2TS \add_x_22_0/U3  (.S(\addr_calc/fft_read_calc/counter/N72 ), 
	.CO(\add_x_22_0/n2 ), 
	.CIN(\add_x_22_0/n3 ), 
	.A(\addr_calc/fft_read_calc/count[29] ));
   DFFHQX2TS \addr_calc/iir_read_calc/counter/count_reg[8]  (.Q(\addr_calc/iir_read_calc/count[8] ), 
	.D(n963), 
	.CK(clk__L1_N0));
   DFFX4TS \addr_calc/fir_read_calc/counter/count_reg[26]  (.Q(\addr_calc/fir_read_calc/count[26] ), 
	.D(n1072), 
	.CK(clk__L1_N0));
   DFFHQX2TS \addr_calc/fir_write_calc/counter/count_reg[26]  (.Q(\addr_calc/fir_write_calc/count[26] ), 
	.D(n1104), 
	.CK(clk__L1_N0));
   DFFHQX4TS \addr_calc/iir_write_calc/counter/count_reg[22]  (.Q(\addr_calc/iir_write_calc/count[22] ), 
	.D(n980), 
	.CK(clk__L1_N0));
   DFFHQX4TS \addr_calc/fir_write_calc/counter/count_reg[24]  (.Q(\addr_calc/fir_write_calc/count[24] ), 
	.D(n1106), 
	.CK(clk__L1_N0));
   DFFHQX4TS \addr_calc/iir_read_calc/counter/count_reg[26]  (.Q(\addr_calc/iir_read_calc/count[26] ), 
	.D(n945), 
	.CK(clk__L1_N0));
   DFFHQX1TS \addr_calc/fft_read_calc/counter/count_reg[26]  (.Q(\addr_calc/fft_read_calc/count[26] ), 
	.D(n1008), 
	.CK(clk__L1_N0));
   DFFHQX4TS \addr_calc/fft_write_calc/counter/count_reg[26]  (.Q(\addr_calc/fft_write_calc/count[26] ), 
	.D(n1040), 
	.CK(clk__L1_N0));
   DFFHQX4TS \addr_calc/iir_write_calc/counter/count_reg[26]  (.Q(\addr_calc/iir_write_calc/count[26] ), 
	.D(n976), 
	.CK(clk__L1_N0));
   DFFQX1TS \addr_calc/iir_write_calc/counter/count_reg[18]  (.Q(\addr_calc/iir_write_calc/count[18] ), 
	.D(n984), 
	.CK(clk__L1_N0));
   DFFHQX1TS \addr_calc/iir_write_calc/counter/count_reg[14]  (.Q(\addr_calc/iir_write_calc/count[14] ), 
	.D(n988), 
	.CK(clk__L1_N0));
   DFFHQX1TS \addr_calc/fft_read_calc/counter/count_reg[18]  (.Q(\addr_calc/fft_read_calc/count[18] ), 
	.D(n1016), 
	.CK(clk__L1_N0));
   DFFHQX8TS \addr_calc/fft_write_calc/counter/count_reg[3]  (.Q(\addr_calc/fft_write_calc/count[3] ), 
	.D(n1063), 
	.CK(clk__L1_N0));
   DFFHQX4TS \addr_calc/fft_write_calc/counter/count_reg[16]  (.Q(\addr_calc/fft_write_calc/count[16] ), 
	.D(n1050), 
	.CK(clk__L1_N0));
   DFFHQX4TS \addr_calc/fir_write_calc/counter/count_reg[16]  (.Q(\addr_calc/fir_write_calc/count[16] ), 
	.D(n1114), 
	.CK(clk__L1_N0));
   DFFHQX4TS \addr_calc/fir_write_calc/counter/count_reg[23]  (.Q(\addr_calc/fir_write_calc/count[23] ), 
	.D(n1107), 
	.CK(clk__L1_N0));
   DFFHQX4TS \addr_calc/iir_write_calc/counter/count_reg[9]  (.Q(\addr_calc/iir_write_calc/count[9] ), 
	.D(n993), 
	.CK(clk__L1_N0));
   DFFHQX4TS \addr_calc/fft_read_calc/counter/count_reg[9]  (.Q(\addr_calc/fft_read_calc/count[9] ), 
	.D(n1025), 
	.CK(clk__L1_N0));
   DFFHQX1TS \addr_calc/fir_read_calc/counter/count_reg[23]  (.Q(\addr_calc/fir_read_calc/count[23] ), 
	.D(n1075), 
	.CK(clk__L1_N0));
   DFFHQX4TS \addr_calc/fft_write_calc/counter/count_reg[28]  (.Q(\addr_calc/fft_write_calc/count[28] ), 
	.D(n1038), 
	.CK(clk__L1_N0));
   DFFHQX4TS \addr_calc/fft_write_calc/counter/count_reg[23]  (.Q(\addr_calc/fft_write_calc/count[23] ), 
	.D(n1043), 
	.CK(clk__L1_N0));
   DFFHQX1TS \addr_calc/fft_read_calc/counter/count_reg[16]  (.Q(\addr_calc/fft_read_calc/count[16] ), 
	.D(n1018), 
	.CK(clk__L1_N0));
   DFFX4TS \addr_calc/fft_read_calc/counter/count_reg[4]  (.Q(\addr_calc/fft_read_calc/count[4] ), 
	.D(n1030), 
	.CK(clk__L1_N0));
   DFFHQX8TS \addr_calc/fir_write_calc/counter/count_reg[31]  (.Q(\addr_calc/fir_write_calc/count[31] ), 
	.D(n1099), 
	.CK(clk__L1_N0));
   DFFHQX2TS \addr_calc/fir_read_calc/counter/count_reg[31]  (.Q(\addr_calc/fir_read_calc/count[31] ), 
	.D(n1132), 
	.CK(clk__L1_N0));
   DFFHQX4TS \addr_calc/fft_read_calc/counter/count_reg[2]  (.Q(\addr_calc/fft_read_calc/count[2] ), 
	.D(n1032), 
	.CK(clk__L1_N0));
   DFFHQX4TS \addr_calc/fft_read_calc/counter/count_reg[8]  (.Q(\addr_calc/fft_read_calc/count[8] ), 
	.D(n1026), 
	.CK(clk__L1_N0));
   DFFHQX8TS \addr_calc/iir_write_calc/counter/count_reg[12]  (.Q(\addr_calc/iir_write_calc/count[12] ), 
	.D(n990), 
	.CK(clk__L1_N0));
   DFFHQX8TS \addr_calc/iir_write_calc/counter/count_reg[8]  (.Q(\addr_calc/iir_write_calc/count[8] ), 
	.D(n994), 
	.CK(clk__L1_N0));
   DFFQX4TS \addr_calc/fft_write_calc/counter/count_reg[0]  (.Q(\addr_calc/fft_write_calc/count[0] ), 
	.D(n1066), 
	.CK(clk__L1_N0));
   DFFHQX8TS \addr_calc/fft_write_calc/counter/count_reg[2]  (.Q(\addr_calc/fft_write_calc/count[2] ), 
	.D(n1064), 
	.CK(clk__L1_N0));
   DFFHQX4TS \addr_calc/fft_write_calc/counter/count_reg[8]  (.Q(\addr_calc/fft_write_calc/count[8] ), 
	.D(n1058), 
	.CK(clk__L1_N0));
   DFFHQX4TS \addr_calc/fft_write_calc/counter/count_reg[12]  (.Q(\addr_calc/fft_write_calc/count[12] ), 
	.D(n1054), 
	.CK(clk__L1_N0));
   DFFQX4TS \addr_calc/fft_write_calc/counter/count_reg[14]  (.Q(\addr_calc/fft_write_calc/count[14] ), 
	.D(n1052), 
	.CK(clk__L1_N0));
   DFFHQX8TS \addr_calc/iir_read_calc/counter/count_reg[6]  (.Q(\addr_calc/iir_read_calc/count[6] ), 
	.D(n965), 
	.CK(clk__L1_N0));
   DFFHQX8TS \addr_calc/iir_read_calc/counter/count_reg[2]  (.Q(\addr_calc/iir_read_calc/count[2] ), 
	.D(n969), 
	.CK(clk__L1_N0));
   DFFHQX4TS \addr_calc/fir_read_calc/counter/count_reg[2]  (.Q(\addr_calc/fir_read_calc/count[2] ), 
	.D(n1096), 
	.CK(clk__L1_N0));
   DFFHQX4TS \addr_calc/fir_read_calc/counter/count_reg[6]  (.Q(\addr_calc/fir_read_calc/count[6] ), 
	.D(n1092), 
	.CK(clk__L1_N0));
   DFFHQX4TS \addr_calc/fir_read_calc/counter/count_reg[8]  (.Q(\addr_calc/fir_read_calc/count[8] ), 
	.D(n1090), 
	.CK(clk__L1_N0));
   DFFQX4TS \addr_calc/fir_write_calc/counter/count_reg[8]  (.Q(\addr_calc/fir_write_calc/count[8] ), 
	.D(n1122), 
	.CK(clk__L1_N0));
   DFFHQX4TS \addr_calc/fir_read_calc/counter/count_reg[12]  (.Q(\addr_calc/fir_read_calc/count[12] ), 
	.D(n1086), 
	.CK(clk__L1_N0));
   DFFHQX8TS \addr_calc/fir_write_calc/counter/count_reg[6]  (.Q(\addr_calc/fir_write_calc/count[6] ), 
	.D(n1124), 
	.CK(clk__L1_N0));
   DFFQX4TS \addr_calc/fir_write_calc/counter/count_reg[0]  (.Q(\addr_calc/fir_write_calc/count[0] ), 
	.D(n1130), 
	.CK(clk__L1_N0));
   DFFHQX4TS \addr_calc/fft_read_calc/counter/count_reg[1]  (.Q(\addr_calc/fft_read_calc/count[1] ), 
	.D(n1033), 
	.CK(clk__L1_N0));
   DFFHQX4TS \addr_calc/fft_read_calc/counter/count_reg[3]  (.Q(\addr_calc/fft_read_calc/count[3] ), 
	.D(n1031), 
	.CK(clk__L1_N0));
   DFFHQX8TS \addr_calc/fft_read_calc/counter/count_reg[5]  (.Q(\addr_calc/fft_read_calc/count[5] ), 
	.D(n1029), 
	.CK(clk__L1_N0));
   DFFHQX4TS \addr_calc/fft_read_calc/counter/count_reg[10]  (.Q(\addr_calc/fft_read_calc/count[10] ), 
	.D(n1024), 
	.CK(clk__L1_N0));
   DFFHQX4TS \addr_calc/fft_read_calc/counter/count_reg[11]  (.Q(\addr_calc/fft_read_calc/count[11] ), 
	.D(n1023), 
	.CK(clk__L1_N0));
   DFFHQX8TS \addr_calc/fft_write_calc/counter/count_reg[1]  (.Q(\addr_calc/fft_write_calc/count[1] ), 
	.D(n1065), 
	.CK(clk__L1_N0));
   DFFHQX8TS \addr_calc/iir_write_calc/counter/count_reg[10]  (.Q(\addr_calc/iir_write_calc/count[10] ), 
	.D(n992), 
	.CK(clk__L1_N0));
   DFFHQX4TS \addr_calc/fft_write_calc/counter/count_reg[7]  (.Q(\addr_calc/fft_write_calc/count[7] ), 
	.D(n1059), 
	.CK(clk__L1_N0));
   DFFHQX8TS \addr_calc/iir_write_calc/counter/count_reg[4]  (.Q(\addr_calc/iir_write_calc/count[4] ), 
	.D(n998), 
	.CK(clk__L1_N0));
   DFFHQX4TS \addr_calc/fft_write_calc/counter/count_reg[9]  (.Q(\addr_calc/fft_write_calc/count[9] ), 
	.D(n1057), 
	.CK(clk__L1_N0));
   DFFQX4TS \addr_calc/iir_write_calc/counter/count_reg[3]  (.Q(\addr_calc/iir_write_calc/count[3] ), 
	.D(n999), 
	.CK(clk__L1_N0));
   DFFHQX4TS \addr_calc/fft_write_calc/counter/count_reg[10]  (.Q(\addr_calc/fft_write_calc/count[10] ), 
	.D(n1056), 
	.CK(clk__L1_N0));
   DFFHQX8TS \addr_calc/iir_write_calc/counter/count_reg[1]  (.Q(\addr_calc/iir_write_calc/count[1] ), 
	.D(n1001), 
	.CK(clk__L1_N0));
   DFFHQX4TS \addr_calc/fft_write_calc/counter/count_reg[17]  (.Q(\addr_calc/fft_write_calc/count[17] ), 
	.D(n1049), 
	.CK(clk__L1_N0));
   DFFQX4TS \addr_calc/fir_read_calc/counter/count_reg[1]  (.Q(\addr_calc/fir_read_calc/count[1] ), 
	.D(n1097), 
	.CK(clk__L1_N0));
   DFFQX4TS \addr_calc/iir_read_calc/counter/count_reg[10]  (.Q(\addr_calc/iir_read_calc/count[10] ), 
	.D(n961), 
	.CK(clk__L1_N0));
   DFFHQX4TS \addr_calc/fir_read_calc/counter/count_reg[3]  (.Q(\addr_calc/fir_read_calc/count[3] ), 
	.D(n1095), 
	.CK(clk__L1_N0));
   DFFHQX4TS \addr_calc/fir_read_calc/counter/count_reg[4]  (.Q(\addr_calc/fir_read_calc/count[4] ), 
	.D(n1094), 
	.CK(clk__L1_N0));
   DFFQX4TS \addr_calc/iir_read_calc/counter/count_reg[7]  (.Q(\addr_calc/iir_read_calc/count[7] ), 
	.D(n964), 
	.CK(clk__L1_N0));
   DFFHQX8TS \addr_calc/fir_read_calc/counter/count_reg[5]  (.Q(\addr_calc/fir_read_calc/count[5] ), 
	.D(n1093), 
	.CK(clk__L1_N0));
   DFFX4TS \addr_calc/iir_read_calc/counter/count_reg[4]  (.Q(\addr_calc/iir_read_calc/count[4] ), 
	.D(n967), 
	.CK(clk__L1_N0));
   DFFHQX8TS \addr_calc/iir_read_calc/counter/count_reg[1]  (.Q(\addr_calc/iir_read_calc/count[1] ), 
	.D(n970), 
	.CK(clk__L1_N0));
   DFFHQX4TS \addr_calc/fir_write_calc/counter/count_reg[28]  (.Q(\addr_calc/fir_write_calc/count[28] ), 
	.D(n1102), 
	.CK(clk__L1_N0));
   DFFHQX4TS \addr_calc/fir_read_calc/counter/count_reg[11]  (.Q(\addr_calc/fir_read_calc/count[11] ), 
	.D(n1087), 
	.CK(clk__L1_N0));
   DFFHQX4TS \addr_calc/fir_read_calc/counter/count_reg[13]  (.Q(\addr_calc/fir_read_calc/count[13] ), 
	.D(n1085), 
	.CK(clk__L1_N0));
   DFFHQX4TS \addr_calc/fir_read_calc/counter/count_reg[15]  (.Q(\addr_calc/fir_read_calc/count[15] ), 
	.D(n1083), 
	.CK(clk__L1_N0));
   DFFHQX4TS \addr_calc/fir_read_calc/counter/count_reg[17]  (.Q(\addr_calc/fir_read_calc/count[17] ), 
	.D(n1081), 
	.CK(clk__L1_N0));
   DFFHQX4TS \addr_calc/fir_read_calc/counter/count_reg[19]  (.Q(\addr_calc/fir_read_calc/count[19] ), 
	.D(n1079), 
	.CK(clk__L1_N0));
   DFFHQX4TS \addr_calc/fir_write_calc/counter/count_reg[13]  (.Q(\addr_calc/fir_write_calc/count[13] ), 
	.D(n1117), 
	.CK(clk__L1_N0));
   DFFHQX4TS \addr_calc/fir_write_calc/counter/count_reg[11]  (.Q(\addr_calc/fir_write_calc/count[11] ), 
	.D(n1119), 
	.CK(clk__L1_N0));
   DFFHQX4TS \addr_calc/fir_write_calc/counter/count_reg[10]  (.Q(\addr_calc/fir_write_calc/count[10] ), 
	.D(n1120), 
	.CK(clk__L1_N0));
   DFFQX4TS \addr_calc/fir_read_calc/counter/count_reg[27]  (.Q(\addr_calc/fir_read_calc/count[27] ), 
	.D(n1071), 
	.CK(clk__L1_N0));
   DFFHQX4TS \addr_calc/fir_write_calc/counter/count_reg[7]  (.Q(\addr_calc/fir_write_calc/count[7] ), 
	.D(n1123), 
	.CK(clk__L1_N0));
   DFFHQX2TS \addr_calc/fir_write_calc/counter/count_reg[1]  (.Q(\addr_calc/fir_write_calc/count[1] ), 
	.D(n1129), 
	.CK(clk__L1_N0));
   DFFHQX4TS \addr_calc/fir_write_calc/counter/count_reg[3]  (.Q(\addr_calc/fir_write_calc/count[3] ), 
	.D(n1127), 
	.CK(clk__L1_N0));
   DFFHQX8TS \addr_calc/fir_write_calc/counter/count_reg[4]  (.Q(\addr_calc/fir_write_calc/count[4] ), 
	.D(n1126), 
	.CK(clk__L1_N0));
   DFFHQX4TS \addr_calc/iir_write_calc/counter/count_reg[31]  (.Q(\addr_calc/iir_write_calc/count[31] ), 
	.D(n1136), 
	.CK(clk__L1_N0));
   DFFHQX4TS \addr_calc/iir_write_calc/counter/count_reg[30]  (.Q(\addr_calc/iir_write_calc/count[30] ), 
	.D(n1003), 
	.CK(clk__L1_N0));
   DFFHQX8TS \addr_calc/fir_write_calc/counter/count_reg[30]  (.Q(\addr_calc/fir_write_calc/count[30] ), 
	.D(n1100), 
	.CK(clk__L1_N0));
   TBUFX4TS \addr_calc/addr_tri6[13]  (.Y(addr[13]), 
	.OE(n3), 
	.A(\addr_calc/iir_write_addr[13] ));
   DFFQX2TS \addr_calc/iir_read_calc/counter/count_reg[12]  (.Q(\addr_calc/iir_read_calc/count[12] ), 
	.D(n959), 
	.CK(clk__L1_N0));
   DFFTRX2TS \addr_calc/fft_read_calc/counter/done_reg  (.RN(n2072), 
	.QN(n895), 
	.Q(fft_read_done), 
	.D(n783), 
	.CK(clk__L1_N0));
   DFFHQX8TS \addr_calc/iir_read_calc/counter/count_reg[28]  (.Q(\addr_calc/iir_read_calc/count[28] ), 
	.D(n943), 
	.CK(clk__L1_N0));
   DFFQX4TS \addr_calc/iir_read_calc/counter/count_reg[11]  (.Q(\addr_calc/iir_read_calc/count[11] ), 
	.D(n960), 
	.CK(clk__L1_N0));
   DFFHQX4TS \addr_calc/iir_read_calc/counter/count_reg[13]  (.Q(\addr_calc/iir_read_calc/count[13] ), 
	.D(n958), 
	.CK(clk__L1_N0));
   TBUFX6TS \addr_calc/addr_tri5[18]  (.Y(addr[18]), 
	.OE(FE_OFN157_n67), 
	.A(\addr_calc/iir_read_addr[18] ));
   DFFTRX2TS \addr_calc/iir_write_calc/counter/done_reg  (.RN(iir_enable), 
	.Q(iir_write_done), 
	.D(n787), 
	.CK(clk__L1_N0));
   DFFHQX2TS \addr_calc/iir_read_calc/counter/count_reg[19]  (.Q(\addr_calc/iir_read_calc/count[19] ), 
	.D(n952), 
	.CK(clk__L1_N0));
   DFFTRX2TS \addr_calc/fir_read_calc/counter/done_reg  (.RN(FE_OFN564_n2066), 
	.QN(n900), 
	.Q(fir_read_done), 
	.D(n1461), 
	.CK(clk__L1_N0));
   DFFQX4TS \addr_calc/iir_read_calc/counter/count_reg[27]  (.Q(\addr_calc/iir_read_calc/count[27] ), 
	.D(n944), 
	.CK(clk__L1_N0));
   DFFQX4TS \addr_calc/iir_read_calc/counter/count_reg[31]  (.Q(\addr_calc/iir_read_calc/count[31] ), 
	.D(n972), 
	.CK(clk__L1_N0));
   DFFQX4TS \addr_calc/fft_read_calc/counter/count_reg[28]  (.Q(\addr_calc/fft_read_calc/count[28] ), 
	.D(n1006), 
	.CK(clk__L1_N0));
   DFFQX4TS \addr_calc/fft_read_calc/counter/count_reg[20]  (.Q(\addr_calc/fft_read_calc/count[20] ), 
	.D(n1014), 
	.CK(clk__L1_N0));
   DFFTRX2TS \addr_calc/fir_write_calc/counter/done_reg  (.RN(fir_enable), 
	.Q(fir_write_done), 
	.D(n785), 
	.CK(clk__L1_N0));
   DFFQX1TS \addr_calc/fir_write_calc/counter/count_reg[12]  (.Q(\addr_calc/fir_write_calc/count[12] ), 
	.D(n1118), 
	.CK(clk__L1_N0));
   DFFQX4TS \addr_calc/fir_write_calc/counter/count_reg[25]  (.Q(\addr_calc/fir_write_calc/count[25] ), 
	.D(n1105), 
	.CK(clk__L1_N0));
   AOI22XLTS U361 (.Y(n930), 
	.B1(FE_OFN516_from_iir_full), 
	.B0(FE_OFN515_from_iir_empty), 
	.A1(FE_OFN514_to_iir_full), 
	.A0(FE_OFN513_to_iir_empty));
   NAND2BXLTS U374 (.Y(n938), 
	.B(FE_OFN508_from_fft_full), 
	.AN(FE_OFN506_to_fft_full));
   NAND2XLTS \add_x_19_3/U5  (.Y(\add_x_19_3/n34 ), 
	.B(FE_OFN339_offset_31_), 
	.A(FE_OFN262_addr_calc_fir_write_calc_count_31_));
   NAND2X1TS \DP_OP_158_296_6262/U1804  (.Y(\DP_OP_158_296_6262/n1829 ), 
	.B(\DP_OP_158_296_6262/n1830 ), 
	.A(\DP_OP_158_296_6262/n1837 ));
   NAND2XLTS \add_x_22_5/U13  (.Y(\add_x_22_5/n10 ), 
	.B(\addr_calc/iir_write_calc/count[27] ), 
	.A(n2573));
   NAND2XLTS \add_x_22_0/U13  (.Y(\add_x_22_0/n10 ), 
	.B(\addr_calc/fft_read_calc/count[27] ), 
	.A(n2575));
   NAND2XLTS \add_x_22_1/U13  (.Y(\add_x_22_1/n10 ), 
	.B(\addr_calc/fft_write_calc/count[27] ), 
	.A(n2574));
   NAND2XLTS \add_x_22_3/U13  (.Y(\add_x_22_3/n10 ), 
	.B(\addr_calc/fir_write_calc/count[27] ), 
	.A(FE_OFN268_addr_calc_fir_write_calc_count_26_));
   NAND2XLTS \add_x_22_2/U13  (.Y(\add_x_22_2/n10 ), 
	.B(FE_OFN243_addr_calc_fir_read_calc_count_27_), 
	.A(FE_OFN270_addr_calc_fir_read_calc_count_26_));
   NOR2X4TS \add_x_19_0/U104  (.Y(\add_x_19_0/n97 ), 
	.B(FE_OCPUNCON1079_FE_OFN382_offset_19_), 
	.A(n1956));
   OAI32X1TS U354 (.Y(n928), 
	.B1(n2073), 
	.B0(FE_OFN564_n2066), 
	.A2(fir_write_done), 
	.A1(n2071), 
	.A0(fir_read_done));
   NAND2XLTS \add_x_19_0/U5  (.Y(\add_x_19_0/n34 ), 
	.B(FE_OFN339_offset_31_), 
	.A(FE_OFN226_addr_calc_fft_read_calc_count_31_));
   OAI21X1TS \add_x_19_5/U239  (.Y(\add_x_19_5/n183 ), 
	.B0(\add_x_19_5/n185 ), 
	.A1(\add_x_19_5/n184 ), 
	.A0(\add_x_19_5/n186 ));
   NOR3X1TS U356 (.Y(n797), 
	.C(FE_OFN561_n2587), 
	.B(fft_read_done), 
	.A(n1478));
   NAND2X2TS \add_x_19_2/U67  (.Y(\add_x_19_2/n74 ), 
	.B(\add_x_19_2/n76 ), 
	.A(\add_x_19_2/n84 ));
   NAND2XLTS \add_x_22_5/U7  (.Y(\add_x_22_5/n5 ), 
	.B(n1974), 
	.A(\add_x_22_5/n9 ));
   NAND3XLTS U367 (.Y(\data_cntl/N255 ), 
	.C(n2585), 
	.B(n934), 
	.A(FE_OFN566_n2066));
   AND2X2TS U389 (.Y(n936), 
	.B(n2585), 
	.A(FE_OFN566_n2066));
   NOR2X4TS \add_x_19_0/U24  (.Y(\add_x_19_0/n46 ), 
	.B(\add_x_19_0/n48 ), 
	.A(\add_x_19_0/n51 ));
   OAI211X1TS U348 (.Y(n926), 
	.C0(n898), 
	.B0(iir_enable), 
	.A1(FE_OFN563_n2060), 
	.A0(n1829));
   CLKINVX1TS U344 (.Y(n923), 
	.A(n792));
   AOI211XLTS U363 (.Y(\data_cntl/N257 ), 
	.C0(n932), 
	.B0(FE_OFN515_from_iir_empty), 
	.A1(n931), 
	.A0(FE_OFN513_to_iir_empty));
   NAND2XLTS \add_x_22_3/U112  (.Y(\add_x_22_3/n90 ), 
	.B(FE_OFN256_addr_calc_fir_write_calc_count_8_), 
	.A(\add_x_22_3/n93 ));
   OR3XLTS U360 (.Y(\data_cntl/N258 ), 
	.C(n930), 
	.B(\data_cntl/N263 ), 
	.A(FE_OFN151_n2074));
   NAND2XLTS \add_x_22_5/U112  (.Y(\add_x_22_5/n90 ), 
	.B(n2041), 
	.A(\add_x_22_5/n93 ));
   NOR2X1TS U392 (.Y(\data_cntl/N259 ), 
	.B(FE_OFN332_data_cntl_N63), 
	.A(n2585));
   NOR3X1TS U393 (.Y(\data_cntl/N261 ), 
	.C(n2585), 
	.B(FE_OFN322_data_cntl_N9), 
	.A(FE_OFN333_data_to_fft));
   NAND3XLTS U395 (.Y(\addr_calc/N216 ), 
	.C(FE_OFN333_data_to_fft), 
	.B(FE_OFN323_data_from_fft), 
	.A(n2071));
   AOI211XLTS U369 (.Y(\data_cntl/N254 ), 
	.C0(n1830), 
	.B0(FE_OFN511_from_fir_empty), 
	.A1(n935), 
	.A0(FE_OFN509_to_fir_empty));
   CLKINVX1TS U305 (.Y(n888), 
	.A(n899));
   CLKINVX2TS U304 (.Y(n887), 
	.A(n870));
   NOR3X1TS U378 (.Y(\data_cntl/N267 ), 
	.C(n932), 
	.B(FE_OFN314_data_cntl_N159), 
	.A(FE_OFN327_data_to_iir));
   NOR2X1TS U380 (.Y(\data_cntl/N265 ), 
	.B(n932), 
	.A(FE_OFN326_data_cntl_N191));
   NAND4X1TS U382 (.Y(\addr_calc/N224 ), 
	.D(n1830), 
	.C(n940), 
	.B(FE_OFN315_data_from_iir), 
	.A(FE_OFN327_data_to_iir));
   AND2X2TS U355 (.Y(fft_put_req), 
	.B(fft_put_req_reg), 
	.A(n797));
   OAI211XLTS U302 (.Y(n890), 
	.C0(acc_done), 
	.B0(n873), 
	.A1(n901), 
	.A0(n888));
   NAND4BXLTS U278 (.Y(n871), 
	.D(n873), 
	.C(n2074), 
	.B(FE_OFN145_n801), 
	.AN(n872));
   NOR2X1TS U388 (.Y(\data_cntl/N262 ), 
	.B(n1830), 
	.A(FE_OFN329_data_cntl_N99));
   NAND4X1TS U390 (.Y(\addr_calc/N220 ), 
	.D(n2588), 
	.C(FE_OFN319_data_from_fir), 
	.B(FE_OFN330_data_to_fir), 
	.A(FE_OFN565_n2066));
   NAND2BXLTS U364 (.Y(n931), 
	.B(FE_OFN516_from_iir_full), 
	.AN(FE_OFN514_to_iir_full));
   NOR2XLTS U366 (.Y(n933), 
	.B(FE_OFN515_from_iir_empty), 
	.A(FE_OFN513_to_iir_empty));
   NAND2BX1TS U370 (.Y(n935), 
	.B(FE_OFN512_from_fir_full), 
	.AN(FE_OFN510_to_fir_full));
   NOR2XLTS U372 (.Y(n937), 
	.B(FE_OFN511_from_fir_empty), 
	.A(FE_OFN509_to_fir_empty));
   AO22X1TS U368 (.Y(n934), 
	.B1(FE_OFN512_from_fir_full), 
	.B0(FE_OFN511_from_fir_empty), 
	.A1(FE_OFN510_to_fir_full), 
	.A0(FE_OFN509_to_fir_empty));
   NOR2X1TS \add_x_19_4/U38  (.Y(\add_x_19_4/n55 ), 
	.B(FE_OFN355_offset_27_), 
	.A(FE_OFN235_addr_calc_iir_read_calc_count_27_));
   NOR3XLTS U375 (.Y(\data_cntl/N251 ), 
	.C(n939), 
	.B(FE_OFN506_to_fft_full), 
	.A(FE_OFN508_from_fft_full));
   NOR2X2TS \add_x_19_2/U69  (.Y(\add_x_19_2/n76 ), 
	.B(\add_x_19_2/n78 ), 
	.A(\add_x_19_2/n81 ));
   NAND2XLTS \add_x_22_5/U143  (.Y(\add_x_22_5/n115 ), 
	.B(n2036), 
	.A(\add_x_22_5/n118 ));
   NAND2X2TS \add_x_19_5/U67  (.Y(\add_x_19_5/n74 ), 
	.B(\add_x_19_5/n76 ), 
	.A(\add_x_19_5/n84 ));
   NAND2X1TS \add_x_22_1/U7  (.Y(\add_x_22_1/n5 ), 
	.B(n2557), 
	.A(\add_x_22_1/n9 ));
   NOR2X2TS \add_x_19_3/U34  (.Y(\add_x_19_3/n53 ), 
	.B(\add_x_19_3/n55 ), 
	.A(\add_x_19_3/n58 ));
   NOR2X2TS \add_x_19_5/U24  (.Y(\add_x_19_5/n46 ), 
	.B(\add_x_19_5/n48 ), 
	.A(\add_x_19_5/n51 ));
   NAND3XLTS U345 (.Y(n792), 
	.C(n924), 
	.B(iir_read_done), 
	.A(n2063));
   NAND2X1TS \add_x_22_2/U123  (.Y(\add_x_22_2/n99 ), 
	.B(n2001), 
	.A(\add_x_22_2/n102 ));
   NOR2X2TS \add_x_19_1/U24  (.Y(\add_x_19_1/n46 ), 
	.B(\add_x_19_1/n48 ), 
	.A(\add_x_19_1/n51 ));
   NAND2X1TS \add_x_22_0/U112  (.Y(\add_x_22_0/n90 ), 
	.B(n2049), 
	.A(\add_x_22_0/n93 ));
   NAND2XLTS U308 (.Y(n901), 
	.B(n884), 
	.A(n870));
   NAND2X1TS \add_x_22_1/U81  (.Y(\add_x_22_1/n65 ), 
	.B(FE_OFN259_addr_calc_fft_write_calc_count_14_), 
	.A(\add_x_22_1/n68 ));
   NAND2X1TS \add_x_22_1/U59  (.Y(\add_x_22_1/n47 ), 
	.B(\addr_calc/fft_write_calc/count[18] ), 
	.A(\add_x_22_1/n50 ));
   NAND2X1TS \add_x_22_1/U39  (.Y(\add_x_22_1/n31 ), 
	.B(FE_OFN285_addr_calc_fft_write_calc_count_22_), 
	.A(\add_x_22_1/n34 ));
   NAND2X1TS \add_x_22_0/U81  (.Y(\add_x_22_0/n65 ), 
	.B(\addr_calc/fft_read_calc/count[14] ), 
	.A(\add_x_22_0/n68 ));
   AND2X2TS U349 (.Y(fir_put_req), 
	.B(fir_put_req_reg), 
	.A(n798));
   NOR2X1TS \add_x_19_1/U178  (.Y(\add_x_19_1/n144 ), 
	.B(FE_OFN418_offset_10_), 
	.A(\addr_calc/fft_write_calc/count[10] ));
   NAND2X1TS \add_x_22_3/U35  (.Y(\add_x_22_3/n28 ), 
	.B(n2563), 
	.A(n1668));
   NOR2X2TS \add_x_19_5/U69  (.Y(\add_x_19_5/n76 ), 
	.B(\add_x_19_5/n78 ), 
	.A(\add_x_19_5/n81 ));
   NAND2X2TS \add_x_19_4/U67  (.Y(\add_x_19_4/n74 ), 
	.B(\add_x_19_4/n76 ), 
	.A(\add_x_19_4/n84 ));
   NOR2XLTS \add_x_22_2/U132  (.Y(\add_x_22_2/n106 ), 
	.B(\add_x_22_2/n109 ), 
	.A(\add_x_22_2/n110 ));
   NAND2XLTS \add_x_22_4/U112  (.Y(\add_x_22_4/n90 ), 
	.B(n2583), 
	.A(\add_x_22_4/n93 ));
   NAND2XLTS \add_x_22_1/U112  (.Y(\add_x_22_1/n90 ), 
	.B(n2026), 
	.A(\add_x_22_1/n93 ));
   NAND2XLTS \add_x_22_2/U112  (.Y(\add_x_22_2/n90 ), 
	.B(n1997), 
	.A(\add_x_22_2/n93 ));
   NAND2XLTS \add_x_22_0/U123  (.Y(\add_x_22_0/n99 ), 
	.B(FE_OFN225_addr_calc_fft_read_calc_count_6_), 
	.A(\add_x_22_0/n102 ));
   DFFHQX4TS \addr_calc/iir_write_calc/counter/count_reg[6]  (.Q(\addr_calc/iir_write_calc/count[6] ), 
	.D(n996), 
	.CK(clk__L1_N0));
   DFFHQX1TS \addr_calc/iir_write_calc/counter/count_reg[20]  (.Q(\addr_calc/iir_write_calc/count[20] ), 
	.D(n982), 
	.CK(clk__L1_N0));
   DFFQX1TS \addr_calc/iir_write_calc/counter/count_reg[15]  (.Q(\addr_calc/iir_write_calc/count[15] ), 
	.D(n987), 
	.CK(clk__L1_N0));
   DFFHQX1TS \addr_calc/iir_write_calc/counter/count_reg[16]  (.Q(\addr_calc/iir_write_calc/count[16] ), 
	.D(n986), 
	.CK(clk__L1_N0));
   DFFQX2TS \addr_calc/iir_write_calc/counter/count_reg[29]  (.Q(\addr_calc/iir_write_calc/count[29] ), 
	.D(n973), 
	.CK(clk__L1_N0));
   TBUFX16TS \addr_calc/addr_tri5[21]  (.Y(addr[21]), 
	.OE(FE_OFN158_n67), 
	.A(\addr_calc/iir_read_addr[21] ));
   TBUFX12TS \addr_calc/addr_tri6[21]  (.Y(addr[21]), 
	.OE(FE_OFN154_n3), 
	.A(FE_OFN123_addr_calc_iir_write_addr_21_));
   TBUFX12TS \addr_calc/addr_tri4[21]  (.Y(addr[21]), 
	.OE(FE_OFN174_n131), 
	.A(\addr_calc/fir_write_addr[21] ));
   TBUFX4TS \addr_calc/addr_tri5[24]  (.Y(addr[24]), 
	.OE(FE_OFN294_n2642), 
	.A(FE_OFN116_addr_calc_iir_read_addr_24_));
   NAND2XLTS \DP_OP_158_296_6262/U1847  (.Y(\DP_OP_158_296_6262/n1861 ), 
	.B(\DP_OP_158_296_6262/n1862 ), 
	.A(FE_OFN112_DP_OP_158_296_6262_n1791));
   NAND2X1TS \add_x_19_4/U26  (.Y(\add_x_19_4/n4 ), 
	.B(\add_x_19_4/n49 ), 
	.A(\add_x_19_4/n195 ));
   NAND2X1TS \add_x_19_4/U50  (.Y(\add_x_19_4/n7 ), 
	.B(\add_x_19_4/n64 ), 
	.A(\add_x_19_4/n198 ));
   NAND2X1TS \add_x_19_4/U22  (.Y(\add_x_19_4/n44 ), 
	.B(\add_x_19_4/n46 ), 
	.A(\add_x_19_4/n72 ));
   OAI21X2TS \add_x_19_4/U25  (.Y(\add_x_19_4/n47 ), 
	.B0(\add_x_19_4/n49 ), 
	.A1(\add_x_19_4/n48 ), 
	.A0(\add_x_19_4/n52 ));
   OAI21X2TS \add_x_19_4/U142  (.Y(\add_x_19_4/n122 ), 
	.B0(\add_x_19_4/n124 ), 
	.A1(\add_x_19_4/n123 ), 
	.A0(\add_x_19_4/n125 ));
   NAND2X1TS \add_x_19_4/U137  (.Y(\add_x_19_4/n17 ), 
	.B(\add_x_19_4/n121 ), 
	.A(\add_x_19_4/n208 ));
   NOR2X1TS \add_x_22_1/U132  (.Y(\add_x_22_1/n106 ), 
	.B(\add_x_22_1/n109 ), 
	.A(\add_x_22_1/n110 ));
   NOR2X1TS \DP_OP_159_297_3515/U941  (.Y(\DP_OP_159_297_3515/n942 ), 
	.B(\DP_OP_159_297_3515/n943 ), 
	.A(\DP_OP_159_297_3515/n957 ));
   NAND2X1TS \DP_OP_158_296_6262/U1874  (.Y(\DP_OP_158_296_6262/n1882 ), 
	.B(\DP_OP_158_296_6262/n1904 ), 
	.A(\DP_OP_158_296_6262/n1883 ));
   OAI21X2TS \add_x_19_0/U136  (.Y(\add_x_19_0/n119 ), 
	.B0(\add_x_19_0/n121 ), 
	.A1(\add_x_19_0/n124 ), 
	.A0(\add_x_19_0/n120 ));
   NAND2X2TS \DP_OP_158_296_6262/U1090  (.Y(\DP_OP_158_296_6262/n1071 ), 
	.B(\DP_OP_158_296_6262/n1174 ), 
	.A(\DP_OP_158_296_6262/n1073 ));
   NOR2X2TS \DP_OP_158_296_6262/U1092  (.Y(\DP_OP_158_296_6262/n1073 ), 
	.B(\DP_OP_158_296_6262/n1132 ), 
	.A(\DP_OP_158_296_6262/n1075 ));
   XNOR2X4TS \DP_OP_158_296_6262/U906  (.Y(\DP_OP_158_296_6262/n899 ), 
	.B(FE_OFN226_addr_calc_fft_read_calc_count_31_), 
	.A(n1778));
   XNOR2X1TS \DP_OP_158_296_6262/U1185  (.Y(\DP_OP_158_296_6262/n1160 ), 
	.B(\addr_calc/fft_read_calc/count[13] ), 
	.A(FE_OFN524_n1659));
   XNOR2X1TS \DP_OP_158_296_6262/U1219  (.Y(\DP_OP_158_296_6262/n1191 ), 
	.B(n1972), 
	.A(n1656));
   XNOR2X1TS \DP_OP_158_296_6262/U1229  (.Y(\DP_OP_158_296_6262/n1200 ), 
	.B(n2560), 
	.A(n1469));
   XNOR2X1TS \DP_OP_158_296_6262/U1239  (.Y(\DP_OP_158_296_6262/n1209 ), 
	.B(n2049), 
	.A(n2598));
   NAND2X1TS \DP_OP_158_296_6262/U1255  (.Y(\DP_OP_158_296_6262/n1223 ), 
	.B(n1599), 
	.A(n1602));
   NAND2X1TS \DP_OP_158_296_6262/U1277  (.Y(\DP_OP_158_296_6262/n1243 ), 
	.B(n1601), 
	.A(n1600));
   NAND2X1TS \DP_OP_158_296_6262/U1295  (.Y(\DP_OP_158_296_6262/n1259 ), 
	.B(n1598), 
	.A(\DP_OP_158_296_6262/n1265 ));
   NOR2X1TS \DP_OP_158_296_6262/U1302  (.Y(\DP_OP_158_296_6262/n1265 ), 
	.B(\DP_OP_158_296_6262/n1269 ), 
	.A(\DP_OP_158_296_6262/n1267 ));
   XNOR2X1TS \DP_OP_158_296_6262/U1304  (.Y(\DP_OP_158_296_6262/n1267 ), 
	.B(n2597), 
	.A(\addr_calc/fft_read_calc/count[1] ));
   XNOR2X1TS \DP_OP_158_296_6262/U1311  (.Y(\DP_OP_158_296_6262/n1269 ), 
	.B(n2058), 
	.A(FE_OFN518_n2372));
   NOR2X1TS \DP_OP_158_296_6262/U1821  (.Y(\DP_OP_158_296_6262/n1842 ), 
	.B(FE_OFN466_filesize_28_), 
	.A(\DP_OP_158_296_6262/n1792 ));
   NAND2X2TS \add_x_19_3/U71  (.Y(\add_x_19_3/n9 ), 
	.B(\add_x_19_3/n79 ), 
	.A(\add_x_19_3/n200 ));
   AOI21X4TS \add_x_19_3/U82  (.Y(\add_x_19_3/n83 ), 
	.B0(\add_x_19_3/n85 ), 
	.A1(\add_x_19_3/n84 ), 
	.A0(\add_x_19_3/n92 ));
   NAND2X1TS \add_x_19_5/U2  (.Y(\add_x_19_5/n1 ), 
	.B(\add_x_19_5/n34 ), 
	.A(n1590));
   NAND2XLTS \add_x_19_5/U5  (.Y(\add_x_19_5/n34 ), 
	.B(FE_OFN340_offset_31_), 
	.A(FE_OFN240_addr_calc_iir_write_calc_count_31_));
   NAND2X2TS \add_x_19_4/U199  (.Y(\add_x_19_4/n158 ), 
	.B(\add_x_19_4/n168 ), 
	.A(\add_x_19_4/n160 ));
   OAI21X2TS \add_x_19_4/U202  (.Y(\add_x_19_4/n161 ), 
	.B0(\add_x_19_4/n163 ), 
	.A1(\add_x_19_4/n166 ), 
	.A0(\add_x_19_4/n162 ));
   OAI21X4TS \add_x_19_4/U216  (.Y(\add_x_19_4/n169 ), 
	.B0(\add_x_19_4/n171 ), 
	.A1(\add_x_19_4/n176 ), 
	.A0(\add_x_19_4/n170 ));
   NAND2X2TS \add_x_19_5/U71  (.Y(\add_x_19_5/n9 ), 
	.B(\add_x_19_5/n79 ), 
	.A(\add_x_19_5/n200 ));
   AOI21X4TS \add_x_19_3/U165  (.Y(\add_x_19_3/n136 ), 
	.B0(\add_x_19_3/n138 ), 
	.A1(\add_x_19_3/n150 ), 
	.A0(\add_x_19_3/n137 ));
   OAI21X2TS \add_x_19_3/U167  (.Y(\add_x_19_3/n138 ), 
	.B0(\add_x_19_3/n140 ), 
	.A1(\add_x_19_3/n145 ), 
	.A0(\add_x_19_3/n139 ));
   XOR2X1TS \add_x_22_5/U42  (.Y(\addr_calc/iir_write_calc/counter/N64 ), 
	.B(n1961), 
	.A(\add_x_22_5/n38 ));
   NAND2X1TS \add_x_22_5/U48  (.Y(\add_x_22_5/n38 ), 
	.B(\addr_calc/iir_write_calc/count[20] ), 
	.A(\add_x_22_5/n41 ));
   NOR2X1TS \DP_OP_159_297_3515/U881  (.Y(\DP_OP_159_297_3515/n900 ), 
	.B(\DP_OP_159_297_3515/n901 ), 
	.A(FE_OFN114_DP_OP_159_297_3515_n852));
   NOR2X1TS \DP_OP_159_297_3515/U883  (.Y(\DP_OP_159_297_3515/n902 ), 
	.B(\DP_OP_159_297_3515/n903 ), 
	.A(\DP_OP_159_297_3515/n915 ));
   NAND2X1TS \DP_OP_159_297_3515/U884  (.Y(\DP_OP_159_297_3515/n903 ), 
	.B(FE_OFN466_filesize_28_), 
	.A(FE_OFN467_filesize_27_));
   NAND2X1TS \DP_OP_159_297_3515/U904  (.Y(\DP_OP_159_297_3515/n915 ), 
	.B(n1664), 
	.A(FE_OFN470_filesize_25_));
   NAND2X2TS \add_x_19_2/U2  (.Y(\add_x_19_2/n1 ), 
	.B(\add_x_19_2/n34 ), 
	.A(n1560));
   NAND2XLTS \add_x_19_2/U5  (.Y(\add_x_19_2/n34 ), 
	.B(FE_OFN337_offset_31_), 
	.A(FE_OFN261_addr_calc_fir_read_calc_count_31_));
   AOI21X4TS \add_x_19_0/U82  (.Y(\add_x_19_0/n83 ), 
	.B0(\add_x_19_0/n85 ), 
	.A1(\add_x_19_0/n84 ), 
	.A0(\add_x_19_0/n92 ));
   OAI21X4TS \add_x_19_0/U97  (.Y(\add_x_19_0/n92 ), 
	.B0(\add_x_19_0/n94 ), 
	.A1(\add_x_19_0/n93 ), 
	.A0(FE_OFN528_add_x_19_0_n113));
   OAI21X1TS \add_x_19_5/U107  (.Y(\add_x_19_5/n99 ), 
	.B0(\add_x_19_5/n101 ), 
	.A1(\add_x_19_5/n100 ), 
	.A0(\add_x_19_5/n102 ));
   NAND2X1TS \add_x_19_5/U102  (.Y(\add_x_19_5/n13 ), 
	.B(\add_x_19_5/n98 ), 
	.A(\add_x_19_5/n204 ));
   NAND2X2TS \add_x_19_1/U36  (.Y(\add_x_19_1/n5 ), 
	.B(\add_x_19_1/n56 ), 
	.A(\add_x_19_1/n196 ));
   NOR2X1TS \add_x_19_1/U232  (.Y(\add_x_19_1/n179 ), 
	.B(\add_x_19_1/n181 ), 
	.A(\add_x_19_1/n184 ));
   OAI21X1TS \add_x_19_1/U233  (.Y(\add_x_19_1/n180 ), 
	.B0(\add_x_19_1/n182 ), 
	.A1(\add_x_19_1/n185 ), 
	.A0(\add_x_19_1/n181 ));
   OAI21X2TS \add_x_19_0/U150  (.Y(\add_x_19_0/n127 ), 
	.B0(\add_x_19_0/n129 ), 
	.A1(\add_x_19_0/n132 ), 
	.A0(\add_x_19_0/n128 ));
   NOR2X2TS \add_x_19_3/U232  (.Y(\add_x_19_3/n179 ), 
	.B(\add_x_19_3/n184 ), 
	.A(\add_x_19_3/n181 ));
   NOR2X8TS \add_x_19_1/U215  (.Y(\add_x_19_1/n168 ), 
	.B(\add_x_19_1/n170 ), 
	.A(\add_x_19_1/n175 ));
   NOR2X8TS \add_x_19_0/U65  (.Y(\add_x_19_0/n72 ), 
	.B(\add_x_19_0/n74 ), 
	.A(\add_x_19_0/n93 ));
   NAND2X4TS \add_x_19_0/U67  (.Y(\add_x_19_0/n74 ), 
	.B(\add_x_19_0/n76 ), 
	.A(\add_x_19_0/n84 ));
   OAI21X4TS \add_x_19_0/U66  (.Y(\add_x_19_0/n73 ), 
	.B0(\add_x_19_0/n75 ), 
	.A1(\add_x_19_0/n74 ), 
	.A0(\add_x_19_0/n94 ));
   AOI21X2TS \add_x_19_0/U68  (.Y(\add_x_19_0/n75 ), 
	.B0(\add_x_19_0/n77 ), 
	.A1(\add_x_19_0/n76 ), 
	.A0(\add_x_19_0/n85 ));
   OAI21X2TS \add_x_19_0/U70  (.Y(\add_x_19_0/n77 ), 
	.B0(\add_x_19_0/n79 ), 
	.A1(\add_x_19_0/n82 ), 
	.A0(\add_x_19_0/n78 ));
   NAND2X1TS \add_x_19_2/U22  (.Y(\add_x_19_2/n44 ), 
	.B(\add_x_19_2/n46 ), 
	.A(\add_x_19_2/n72 ));
   OAI21X2TS \add_x_19_2/U25  (.Y(\add_x_19_2/n47 ), 
	.B0(\add_x_19_2/n49 ), 
	.A1(\add_x_19_2/n48 ), 
	.A0(\add_x_19_2/n52 ));
   NOR2X2TS \add_x_19_0/U135  (.Y(\add_x_19_0/n118 ), 
	.B(\add_x_19_0/n120 ), 
	.A(\add_x_19_0/n123 ));
   NOR2X2TS \add_x_19_1/U166  (.Y(\add_x_19_1/n137 ), 
	.B(\add_x_19_1/n139 ), 
	.A(\add_x_19_1/n144 ));
   NOR2X2TS \add_x_19_1/U135  (.Y(\add_x_19_1/n118 ), 
	.B(\add_x_19_1/n120 ), 
	.A(\add_x_19_1/n123 ));
   NOR2X2TS \add_x_19_2/U24  (.Y(\add_x_19_2/n46 ), 
	.B(\add_x_19_2/n48 ), 
	.A(\add_x_19_2/n51 ));
   NOR2X6TS \add_x_19_1/U201  (.Y(\add_x_19_1/n160 ), 
	.B(\add_x_19_1/n165 ), 
	.A(\add_x_19_1/n162 ));
   OAI21X2TS \add_x_19_2/U216  (.Y(\add_x_19_2/n169 ), 
	.B0(\add_x_19_2/n171 ), 
	.A1(\add_x_19_2/n176 ), 
	.A0(\add_x_19_2/n170 ));
   OAI21X2TS \add_x_19_2/U66  (.Y(\add_x_19_2/n73 ), 
	.B0(\add_x_19_2/n75 ), 
	.A1(\add_x_19_2/n74 ), 
	.A0(\add_x_19_2/n94 ));
   AOI21X2TS \add_x_19_2/U68  (.Y(\add_x_19_2/n75 ), 
	.B0(\add_x_19_2/n77 ), 
	.A1(\add_x_19_2/n85 ), 
	.A0(\add_x_19_2/n76 ));
   OAI21X1TS \add_x_19_2/U70  (.Y(\add_x_19_2/n77 ), 
	.B0(\add_x_19_2/n79 ), 
	.A1(\add_x_19_2/n82 ), 
	.A0(\add_x_19_2/n78 ));
   OAI21X2TS \add_x_19_2/U84  (.Y(\add_x_19_2/n85 ), 
	.B0(\add_x_19_2/n87 ), 
	.A1(\add_x_19_2/n90 ), 
	.A0(\add_x_19_2/n86 ));
   AOI21X4TS \add_x_19_5/U148  (.Y(\add_x_19_5/n125 ), 
	.B0(\add_x_19_5/n127 ), 
	.A1(\add_x_19_5/n126 ), 
	.A0(\add_x_19_5/n134 ));
   OAI21X2TS \add_x_19_5/U25  (.Y(\add_x_19_5/n47 ), 
	.B0(\add_x_19_5/n49 ), 
	.A1(\add_x_19_5/n48 ), 
	.A0(\add_x_19_5/n52 ));
   AOI21X1TS \add_x_19_5/U68  (.Y(\add_x_19_5/n75 ), 
	.B0(\add_x_19_5/n77 ), 
	.A1(\add_x_19_5/n85 ), 
	.A0(\add_x_19_5/n76 ));
   OAI21X2TS \add_x_19_5/U70  (.Y(\add_x_19_5/n77 ), 
	.B0(\add_x_19_5/n79 ), 
	.A1(\add_x_19_5/n82 ), 
	.A0(\add_x_19_5/n78 ));
   OAI21X2TS \add_x_19_5/U84  (.Y(\add_x_19_5/n85 ), 
	.B0(\add_x_19_5/n87 ), 
	.A1(\add_x_19_5/n90 ), 
	.A0(\add_x_19_5/n86 ));
   NAND2X1TS \add_x_19_1/U71  (.Y(\add_x_19_1/n9 ), 
	.B(\add_x_19_1/n79 ), 
	.A(\add_x_19_1/n200 ));
   DFFTRX2TS \addr_calc/fft_write_calc/counter/done_reg  (.RN(n2072), 
	.QN(n1828), 
	.Q(n1478), 
	.D(n1675), 
	.CK(clk__L1_N0));
   DFFTRX2TS \addr_calc/iir_read_calc/counter/done_reg  (.RN(n2063), 
	.QN(n898), 
	.Q(iir_read_done), 
	.D(n1781), 
	.CK(clk__L1_N0));
   DFFXLTS \pla_top/fft_enable_reg  (.QN(n2070), 
	.Q(FE_OFN228_fft_enable), 
	.D(n1131), 
	.CK(clk__L1_N0));
   DFFQX4TS \addr_calc/iir_read_calc/counter/count_reg[14]  (.Q(\addr_calc/iir_read_calc/count[14] ), 
	.D(n957), 
	.CK(clk__L1_N0));
   TBUFX16TS \addr_calc/addr_tri[22]  (.Y(addr[22]), 
	.OE(FE_OFN162_n323), 
	.A(\addr_calc/fft_read_addr[22] ));
   TBUFX8TS \addr_calc/addr_tri6[22]  (.Y(addr[22]), 
	.OE(FE_OFN154_n3), 
	.A(\addr_calc/iir_write_addr[22] ));
   DFFHQX8TS \addr_calc/fir_read_calc/counter/count_reg[7]  (.Q(\addr_calc/fir_read_calc/count[7] ), 
	.D(n1091), 
	.CK(clk__L1_N0));
   DFFHQX8TS \addr_calc/fft_read_calc/counter/count_reg[31]  (.Q(\addr_calc/fft_read_calc/count[31] ), 
	.D(n1035), 
	.CK(clk__L1_N0));
   DFFHQX4TS \addr_calc/fft_read_calc/counter/count_reg[23]  (.Q(\addr_calc/fft_read_calc/count[23] ), 
	.D(n1011), 
	.CK(clk__L1_N0));
   DFFHQX4TS \addr_calc/iir_write_calc/counter/count_reg[23]  (.Q(\addr_calc/iir_write_calc/count[23] ), 
	.D(n979), 
	.CK(clk__L1_N0));
   DFFHQX4TS \addr_calc/iir_write_calc/counter/count_reg[24]  (.Q(\addr_calc/iir_write_calc/count[24] ), 
	.D(n978), 
	.CK(clk__L1_N0));
   TBUFX12TS \addr_calc/addr_tri5[19]  (.Y(addr[19]), 
	.OE(FE_OFN157_n67), 
	.A(\addr_calc/iir_read_addr[19] ));
   TBUFX16TS \addr_calc/addr_tri6[19]  (.Y(addr[19]), 
	.OE(FE_OFN153_n3), 
	.A(FE_OFN125_addr_calc_iir_write_addr_19_));
   TBUFX16TS \addr_calc/addr_tri4[19]  (.Y(addr[19]), 
	.OE(FE_OFN173_n131), 
	.A(\addr_calc/fir_write_addr[19] ));
   TBUFX8TS \addr_calc/addr_tri3[18]  (.Y(addr[18]), 
	.OE(FE_OFN169_n195), 
	.A(\addr_calc/fir_read_addr[18] ));
   DFFHQX4TS \addr_calc/iir_read_calc/counter/count_reg[17]  (.Q(\addr_calc/iir_read_calc/count[17] ), 
	.D(n954), 
	.CK(clk__L1_N0));
   TBUFX4TS \addr_calc/addr_tri6[18]  (.Y(addr[18]), 
	.OE(FE_OFN153_n3), 
	.A(\addr_calc/iir_write_addr[18] ));
   TBUFX4TS \addr_calc/addr_tri2[18]  (.Y(addr[18]), 
	.OE(FE_OFN165_n259), 
	.A(\addr_calc/fft_write_addr[18] ));
   TBUFX16TS \addr_calc/addr_tri4[13]  (.Y(addr[13]), 
	.OE(n131), 
	.A(\addr_calc/fir_write_addr[13] ));
   TBUFX8TS \addr_calc/addr_tri2[13]  (.Y(addr[13]), 
	.OE(n259), 
	.A(\addr_calc/fft_write_addr[13] ));
   TBUFX12TS \addr_calc/addr_tri2[30]  (.Y(addr[30]), 
	.OE(FE_OFN304_n2645), 
	.A(\addr_calc/fft_write_addr[30] ));
   DFFHQX8TS \addr_calc/iir_read_calc/counter/count_reg[23]  (.Q(\addr_calc/iir_read_calc/count[23] ), 
	.D(n948), 
	.CK(clk__L1_N0));
   DFFQX4TS \addr_calc/iir_read_calc/counter/count_reg[15]  (.Q(\addr_calc/iir_read_calc/count[15] ), 
	.D(n956), 
	.CK(clk__L1_N0));
   TBUFX16TS \addr_calc/addr_tri5[25]  (.Y(addr[25]), 
	.OE(FE_OFN295_n2642), 
	.A(\addr_calc/iir_read_addr[25] ));
   TBUFX12TS \addr_calc/addr_tri[25]  (.Y(addr[25]), 
	.OE(FE_OFN299_n2646), 
	.A(\addr_calc/fft_read_addr[25] ));
   TBUFX20TS \addr_calc/addr_tri[28]  (.Y(addr[28]), 
	.OE(FE_OFN298_n2646), 
	.A(FE_OFN133_addr_calc_fft_read_addr_28_));
   TBUFX16TS \addr_calc/addr_tri5[28]  (.Y(addr[28]), 
	.OE(FE_OFN294_n2642), 
	.A(\addr_calc/iir_read_addr[28] ));
   TBUFX16TS \addr_calc/addr_tri2[28]  (.Y(addr[28]), 
	.OE(FE_OFN302_n2645), 
	.A(\addr_calc/fft_write_addr[28] ));
   TBUFX4TS \addr_calc/addr_tri2[14]  (.Y(addr[14]), 
	.OE(n259), 
	.A(\addr_calc/fft_write_addr[14] ));
   TBUFX4TS \addr_calc/addr_tri2[17]  (.Y(addr[17]), 
	.OE(FE_OFN164_n259), 
	.A(\addr_calc/fft_write_addr[17] ));
   TBUFX12TS \addr_calc/addr_tri2[26]  (.Y(addr[26]), 
	.OE(FE_OFN303_n2645), 
	.A(\addr_calc/fft_write_addr[26] ));
   TBUFX12TS \addr_calc/addr_tri2[15]  (.Y(addr[15]), 
	.OE(FE_OFN164_n259), 
	.A(\addr_calc/fft_write_addr[15] ));
   DFFHQX2TS \addr_calc/iir_read_calc/counter/count_reg[22]  (.Q(\addr_calc/iir_read_calc/count[22] ), 
	.D(n949), 
	.CK(clk__L1_N0));
   TBUFX16TS \addr_calc/addr_tri3[21]  (.Y(addr[21]), 
	.OE(FE_OFN170_n195), 
	.A(\addr_calc/fir_read_addr[21] ));
   TBUFX12TS \addr_calc/addr_tri[14]  (.Y(addr[14]), 
	.OE(n323), 
	.A(\addr_calc/fft_read_addr[14] ));
   TBUFX8TS \addr_calc/addr_tri6[30]  (.Y(addr[30]), 
	.OE(FE_OFN292_n2641), 
	.A(\addr_calc/iir_write_addr[30] ));
   TBUFX16TS \addr_calc/addr_tri4[27]  (.Y(addr[27]), 
	.OE(FE_OFN311_n2643), 
	.A(\addr_calc/fir_write_addr[27] ));
   DFFHQX4TS \addr_calc/iir_write_calc/counter/count_reg[2]  (.Q(\addr_calc/iir_write_calc/count[2] ), 
	.D(n1000), 
	.CK(clk__L1_N0));
   DFFHQX4TS \addr_calc/iir_write_calc/counter/count_reg[13]  (.Q(\addr_calc/iir_write_calc/count[13] ), 
	.D(n989), 
	.CK(clk__L1_N0));
   TBUFX8TS \addr_calc/addr_tri5[17]  (.Y(addr[17]), 
	.OE(FE_OFN156_n67), 
	.A(\addr_calc/iir_read_addr[17] ));
   TBUFX12TS \addr_calc/addr_tri5[22]  (.Y(addr[22]), 
	.OE(FE_OFN158_n67), 
	.A(\addr_calc/iir_read_addr[22] ));
   TBUFX16TS \addr_calc/addr_tri3[22]  (.Y(addr[22]), 
	.OE(FE_OFN170_n195), 
	.A(\addr_calc/fir_read_addr[22] ));
   TBUFX12TS \addr_calc/addr_tri2[21]  (.Y(addr[21]), 
	.OE(FE_OFN166_n259), 
	.A(\addr_calc/fft_write_addr[21] ));
   TBUFX16TS \addr_calc/addr_tri[18]  (.Y(addr[18]), 
	.OE(FE_OFN161_n323), 
	.A(\addr_calc/fft_read_addr[18] ));
   TBUFX12TS \addr_calc/addr_tri4[18]  (.Y(addr[18]), 
	.OE(FE_OFN173_n131), 
	.A(\addr_calc/fir_write_addr[18] ));
   TBUFX16TS \addr_calc/addr_tri[23]  (.Y(addr[23]), 
	.OE(FE_OFN162_n323), 
	.A(\addr_calc/fft_read_addr[23] ));
   TBUFX16TS \addr_calc/addr_tri3[23]  (.Y(addr[23]), 
	.OE(FE_OFN170_n195), 
	.A(\addr_calc/fir_read_addr[23] ));
   TBUFX16TS \addr_calc/addr_tri6[23]  (.Y(addr[23]), 
	.OE(FE_OFN154_n3), 
	.A(\addr_calc/iir_write_addr[23] ));
   XOR2X1TS \add_x_22_4/U42  (.Y(\addr_calc/iir_read_calc/counter/N64 ), 
	.B(n1923), 
	.A(\add_x_22_4/n38 ));
   NAND2X1TS \add_x_22_4/U48  (.Y(\add_x_22_4/n38 ), 
	.B(\addr_calc/iir_read_calc/count[20] ), 
	.A(\add_x_22_4/n41 ));
   XNOR2X1TS \DP_OP_159_297_3515/U341  (.Y(\DP_OP_159_297_3515/n312 ), 
	.B(FE_OFN246_addr_calc_iir_read_calc_count_7_), 
	.A(n2609));
   NAND2X1TS \DP_OP_159_297_3515/U347  (.Y(\DP_OP_159_297_3515/n317 ), 
	.B(n1249), 
	.A(n1247));
   NAND2X1TS \DP_OP_159_297_3515/U377  (.Y(\DP_OP_159_297_3515/n343 ), 
	.B(n1246), 
	.A(\DP_OP_159_297_3515/n349 ));
   XNOR2X1TS \DP_OP_159_297_3515/U374  (.Y(\DP_OP_159_297_3515/n341 ), 
	.B(n1902), 
	.A(n2611));
   NOR2X1TS \DP_OP_159_297_3515/U384  (.Y(\DP_OP_159_297_3515/n349 ), 
	.B(\DP_OP_159_297_3515/n353 ), 
	.A(\DP_OP_159_297_3515/n351 ));
   XNOR2X1TS \DP_OP_159_297_3515/U386  (.Y(\DP_OP_159_297_3515/n351 ), 
	.B(\addr_calc/iir_read_calc/count[1] ), 
	.A(FE_OFN501_filesize_1_));
   NAND2X1TS \DP_OP_159_297_3515/U1003  (.Y(\DP_OP_159_297_3515/n986 ), 
	.B(FE_OFN481_filesize_16_), 
	.A(FE_OFN484_filesize_15_));
   XOR2X1TS \add_x_22_3/U115  (.Y(\addr_calc/fir_write_calc/counter/N50 ), 
	.B(\add_x_22_3/n98 ), 
	.A(\add_x_22_3/n99 ));
   NAND2XLTS \add_x_22_3/U123  (.Y(\add_x_22_3/n99 ), 
	.B(FE_OFN254_addr_calc_fir_write_calc_count_6_), 
	.A(\add_x_22_3/n102 ));
   XOR2X1TS \add_x_22_3/U100  (.Y(\addr_calc/fir_write_calc/counter/N53 ), 
	.B(\add_x_22_3/n84 ), 
	.A(\add_x_22_3/n85 ));
   XNOR2X1TS \DP_OP_158_296_6262/U1354  (.Y(\DP_OP_158_296_6262/n1346 ), 
	.B(FE_OFN262_addr_calc_fir_write_calc_count_31_), 
	.A(n1778));
   NOR2X2TS \DP_OP_158_296_6262/U1723  (.Y(\DP_OP_158_296_6262/n1688 ), 
	.B(\DP_OP_158_296_6262/n1706 ), 
	.A(\DP_OP_158_296_6262/n1690 ));
   XNOR2X4TS \DP_OP_158_296_6262/U1406  (.Y(\DP_OP_158_296_6262/n1395 ), 
	.B(\addr_calc/fir_write_calc/count[28] ), 
	.A(n1775));
   XNOR2X1TS \DP_OP_158_296_6262/U1594  (.Y(\DP_OP_158_296_6262/n1571 ), 
	.B(n2564), 
	.A(n2594));
   XNOR2X1TS \DP_OP_158_296_6262/U1621  (.Y(\DP_OP_158_296_6262/n1596 ), 
	.B(n2003), 
	.A(n1657));
   XNOR2X1TS \DP_OP_158_296_6262/U1607  (.Y(\DP_OP_158_296_6262/n1583 ), 
	.B(\addr_calc/fir_write_calc/count[15] ), 
	.A(n1658));
   XNOR2X1TS \DP_OP_158_296_6262/U1655  (.Y(\DP_OP_158_296_6262/n1627 ), 
	.B(n1877), 
	.A(n1660));
   XNOR2X1TS \DP_OP_158_296_6262/U1687  (.Y(\DP_OP_158_296_6262/n1656 ), 
	.B(FE_OFN257_addr_calc_fir_write_calc_count_8_), 
	.A(n2598));
   XNOR2X1TS \DP_OP_158_296_6262/U1695  (.Y(\DP_OP_158_296_6262/n1663 ), 
	.B(n1869), 
	.A(n1651));
   NAND2X2TS \DP_OP_158_296_6262/U1703  (.Y(\DP_OP_158_296_6262/n1670 ), 
	.B(n1236), 
	.A(n1239));
   NAND2X1TS \DP_OP_158_296_6262/U1725  (.Y(\DP_OP_158_296_6262/n1690 ), 
	.B(n1238), 
	.A(n1237));
   NAND2X1TS \DP_OP_158_296_6262/U1743  (.Y(\DP_OP_158_296_6262/n1706 ), 
	.B(n1235), 
	.A(\DP_OP_158_296_6262/n1712 ));
   NOR2X1TS \DP_OP_158_296_6262/U1750  (.Y(\DP_OP_158_296_6262/n1712 ), 
	.B(\DP_OP_158_296_6262/n1716 ), 
	.A(\DP_OP_158_296_6262/n1714 ));
   XNOR2X1TS \DP_OP_158_296_6262/U1752  (.Y(\DP_OP_158_296_6262/n1714 ), 
	.B(FE_OFN242_addr_calc_fir_write_calc_count_1_), 
	.A(n2597));
   NOR2X8TS \DP_OP_158_296_6262/U2008  (.Y(\DP_OP_158_296_6262/n1986 ), 
	.B(\DP_OP_158_296_6262/n1987 ), 
	.A(\DP_OP_158_296_6262/n2011 ));
   XNOR2X1TS \add_x_22_1/U58  (.Y(\addr_calc/fft_write_calc/counter/N61 ), 
	.B(n2019), 
	.A(\add_x_22_1/n50 ));
   NOR2X1TS \DP_OP_158_296_6262/U644  (.Y(\DP_OP_158_296_6262/n626 ), 
	.B(\DP_OP_158_296_6262/n685 ), 
	.A(\DP_OP_158_296_6262/n628 ));
   NOR2X1TS \DP_OP_158_296_6262/U753  (.Y(\DP_OP_158_296_6262/n727 ), 
	.B(FE_OFN540_DP_OP_158_296_6262_n765), 
	.A(\DP_OP_158_296_6262/n729 ));
   NAND2X1TS \DP_OP_158_296_6262/U795  (.Y(\DP_OP_158_296_6262/n765 ), 
	.B(\DP_OP_158_296_6262/n794 ), 
	.A(\DP_OP_158_296_6262/n767 ));
   XNOR2X1TS \DP_OP_158_296_6262/U458  (.Y(\DP_OP_158_296_6262/n452 ), 
	.B(FE_OFN274_addr_calc_fft_write_calc_count_31_), 
	.A(n1778));
   NOR2X1TS \DP_OP_158_296_6262/U827  (.Y(\DP_OP_158_296_6262/n794 ), 
	.B(\DP_OP_158_296_6262/n812 ), 
	.A(\DP_OP_158_296_6262/n796 ));
   XNOR2X1TS \DP_OP_158_296_6262/U698  (.Y(\DP_OP_158_296_6262/n677 ), 
	.B(n2567), 
	.A(n2594));
   XNOR2X1TS \DP_OP_158_296_6262/U737  (.Y(\DP_OP_158_296_6262/n713 ), 
	.B(FE_OFN524_n1659), 
	.A(n1927));
   XNOR2X1TS \DP_OP_158_296_6262/U771  (.Y(\DP_OP_158_296_6262/n744 ), 
	.B(n1932), 
	.A(n1656));
   XNOR2X1TS \DP_OP_158_296_6262/U781  (.Y(\DP_OP_158_296_6262/n753 ), 
	.B(n1934), 
	.A(n1469));
   XNOR2X1TS \DP_OP_158_296_6262/U791  (.Y(\DP_OP_158_296_6262/n762 ), 
	.B(n2026), 
	.A(n2598));
   XNOR2X1TS \DP_OP_158_296_6262/U799  (.Y(\DP_OP_158_296_6262/n769 ), 
	.B(n1936), 
	.A(n1651));
   NAND2X1TS \DP_OP_158_296_6262/U807  (.Y(\DP_OP_158_296_6262/n776 ), 
	.B(n1209), 
	.A(n1212));
   NAND2X1TS \DP_OP_158_296_6262/U829  (.Y(\DP_OP_158_296_6262/n796 ), 
	.B(n1211), 
	.A(n1210));
   NAND2X1TS \DP_OP_158_296_6262/U847  (.Y(\DP_OP_158_296_6262/n812 ), 
	.B(n1208), 
	.A(\DP_OP_158_296_6262/n818 ));
   XNOR2X1TS \DP_OP_158_296_6262/U510  (.Y(\DP_OP_158_296_6262/n501 ), 
	.B(\addr_calc/fft_write_calc/count[28] ), 
	.A(n1775));
   NOR2X1TS \DP_OP_158_296_6262/U854  (.Y(\DP_OP_158_296_6262/n818 ), 
	.B(\DP_OP_158_296_6262/n822 ), 
	.A(\DP_OP_158_296_6262/n820 ));
   XNOR2X1TS \DP_OP_158_296_6262/U856  (.Y(\DP_OP_158_296_6262/n820 ), 
	.B(n1941), 
	.A(n2597));
   NAND2X1TS \DP_OP_158_296_6262/U1883  (.Y(\DP_OP_158_296_6262/n1889 ), 
	.B(\DP_OP_158_296_6262/n1890 ), 
	.A(\DP_OP_158_296_6262/n1904 ));
   XOR2X1TS \add_x_22_4/U131  (.Y(\addr_calc/iir_read_calc/counter/N47 ), 
	.B(\add_x_22_4/n109 ), 
	.A(\add_x_22_4/n110 ));
   XNOR2X1TS \add_x_22_4/U122  (.Y(\addr_calc/iir_read_calc/counter/N49 ), 
	.B(\add_x_22_4/n101 ), 
	.A(\add_x_22_4/n102 ));
   XOR2X1TS \add_x_22_3/U72  (.Y(\addr_calc/fir_write_calc/counter/N58 ), 
	.B(n1882), 
	.A(\add_x_22_3/n65 ));
   OAI21X4TS \add_x_19_2/U31  (.Y(\add_x_19_2/n50 ), 
	.B0(\add_x_19_2/n52 ), 
	.A1(\add_x_19_2/n51 ), 
	.A0(\add_x_19_2/n68 ));
   NAND2X2TS \add_x_19_2/U26  (.Y(\add_x_19_2/n4 ), 
	.B(\add_x_19_2/n49 ), 
	.A(\add_x_19_2/n195 ));
   OAI21X1TS \add_x_19_2/U55  (.Y(\add_x_19_2/n65 ), 
	.B0(\add_x_19_2/n67 ), 
	.A1(\add_x_19_2/n66 ), 
	.A0(\add_x_19_2/n68 ));
   NAND2X1TS \add_x_19_2/U50  (.Y(\add_x_19_2/n7 ), 
	.B(\add_x_19_2/n64 ), 
	.A(\add_x_19_2/n198 ));
   NOR2X2TS \add_x_19_2/U131  (.Y(\add_x_19_2/n114 ), 
	.B(\add_x_19_2/n116 ), 
	.A(\add_x_19_2/n135 ));
   AOI21X2TS \add_x_19_2/U134  (.Y(\add_x_19_2/n117 ), 
	.B0(\add_x_19_2/n119 ), 
	.A1(\add_x_19_2/n127 ), 
	.A0(\add_x_19_2/n118 ));
   OAI21X1TS \add_x_19_2/U136  (.Y(\add_x_19_2/n119 ), 
	.B0(\add_x_19_2/n121 ), 
	.A1(\add_x_19_2/n124 ), 
	.A0(\add_x_19_2/n120 ));
   XOR2X1TS \add_x_22_2/U72  (.Y(\addr_calc/fir_read_calc/counter/N58 ), 
	.B(\add_x_22_2/n64 ), 
	.A(\add_x_22_2/n65 ));
   NAND2X1TS \add_x_22_2/U81  (.Y(\add_x_22_2/n65 ), 
	.B(n1690), 
	.A(\add_x_22_2/n68 ));
   XNOR2X1TS \add_x_22_5/U47  (.Y(\addr_calc/iir_write_calc/counter/N63 ), 
	.B(n2047), 
	.A(\add_x_22_5/n41 ));
   NAND2X1TS \add_x_19_1/U102  (.Y(\add_x_19_1/n13 ), 
	.B(\add_x_19_1/n98 ), 
	.A(\add_x_19_1/n204 ));
   XNOR2X1TS \add_x_22_1/U16  (.Y(\addr_calc/fft_write_calc/counter/N69 ), 
	.B(\add_x_22_1/n15 ), 
	.A(\add_x_22_1/n16 ));
   NOR2X2TS \add_x_19_1/U131  (.Y(\add_x_19_1/n114 ), 
	.B(\add_x_19_1/n116 ), 
	.A(\add_x_19_1/n135 ));
   OAI21X2TS \add_x_19_1/U132  (.Y(\add_x_19_1/n115 ), 
	.B0(\add_x_19_1/n117 ), 
	.A1(\add_x_19_1/n116 ), 
	.A0(\add_x_19_1/n136 ));
   AOI21X1TS \add_x_19_1/U134  (.Y(\add_x_19_1/n117 ), 
	.B0(\add_x_19_1/n119 ), 
	.A1(\add_x_19_1/n127 ), 
	.A0(\add_x_19_1/n118 ));
   OAI21X1TS \add_x_19_1/U136  (.Y(\add_x_19_1/n119 ), 
	.B0(\add_x_19_1/n121 ), 
	.A1(\add_x_19_1/n124 ), 
	.A0(\add_x_19_1/n120 ));
   OAI21X2TS \add_x_19_1/U202  (.Y(\add_x_19_1/n161 ), 
	.B0(\add_x_19_1/n163 ), 
	.A1(\add_x_19_1/n166 ), 
	.A0(\add_x_19_1/n162 ));
   XNOR2X1TS \add_x_22_1/U126  (.Y(\addr_calc/fft_write_calc/counter/N48 ), 
	.B(n1158), 
	.A(\add_x_22_1/n106 ));
   NAND2X1TS \add_x_19_1/U217  (.Y(\add_x_19_1/n27 ), 
	.B(\add_x_19_1/n171 ), 
	.A(\add_x_19_1/n218 ));
   TBUFX8TS \addr_calc/addr_tri3[15]  (.Y(addr[15]), 
	.OE(FE_OFN168_n195), 
	.A(\addr_calc/fir_read_addr[15] ));
   TBUFX20TS \addr_calc/addr_tri[19]  (.Y(addr[19]), 
	.OE(FE_OFN161_n323), 
	.A(\addr_calc/fft_read_addr[19] ));
   DFFHQX1TS \addr_calc/fir_read_calc/counter/count_reg[21]  (.Q(\addr_calc/fir_read_calc/count[21] ), 
	.D(n1077), 
	.CK(clk__L1_N0));
   TBUFX12TS \addr_calc/addr_tri5[15]  (.Y(addr[15]), 
	.OE(FE_OFN156_n67), 
	.A(FE_OFN118_addr_calc_iir_read_addr_15_));
   TBUFX16TS \addr_calc/addr_tri4[28]  (.Y(addr[28]), 
	.OE(FE_OFN310_n2643), 
	.A(\addr_calc/fir_write_addr[28] ));
   DFFHQX4TS \addr_calc/fft_write_calc/counter/count_reg[5]  (.Q(\addr_calc/fft_write_calc/count[5] ), 
	.D(n1061), 
	.CK(clk__L1_N0));
   TBUFX16TS \addr_calc/addr_tri3[25]  (.Y(addr[25]), 
	.OE(FE_OFN307_n2644), 
	.A(\addr_calc/fir_read_addr[25] ));
   TBUFX8TS \addr_calc/addr_tri2[22]  (.Y(addr[22]), 
	.OE(FE_OFN166_n259), 
	.A(\addr_calc/fft_write_addr[22] ));
   TBUFX16TS \addr_calc/addr_tri5[13]  (.Y(addr[13]), 
	.OE(n67), 
	.A(\addr_calc/iir_read_addr[13] ));
   TBUFX4TS \addr_calc/addr_tri3[13]  (.Y(addr[13]), 
	.OE(n195), 
	.A(\addr_calc/fir_read_addr[13] ));
   TBUFX12TS \addr_calc/addr_tri3[28]  (.Y(addr[28]), 
	.OE(FE_OFN306_n2644), 
	.A(\addr_calc/fir_read_addr[28] ));
   TBUFX16TS \addr_calc/addr_tri5[23]  (.Y(addr[23]), 
	.OE(FE_OFN158_n67), 
	.A(\addr_calc/iir_read_addr[23] ));
   TBUFX16TS \addr_calc/addr_tri[15]  (.Y(addr[15]), 
	.OE(FE_OFN160_n323), 
	.A(\addr_calc/fft_read_addr[15] ));
   DFFHQX4TS \addr_calc/iir_write_calc/counter/count_reg[11]  (.Q(\addr_calc/iir_write_calc/count[11] ), 
	.D(n991), 
	.CK(clk__L1_N0));
   TBUFX12TS \addr_calc/addr_tri2[19]  (.Y(addr[19]), 
	.OE(FE_OFN165_n259), 
	.A(\addr_calc/fft_write_addr[19] ));
   TBUFX16TS \addr_calc/addr_tri3[19]  (.Y(addr[19]), 
	.OE(FE_OFN169_n195), 
	.A(\addr_calc/fir_read_addr[19] ));
   TBUFX16TS \addr_calc/addr_tri4[25]  (.Y(addr[25]), 
	.OE(FE_OFN311_n2643), 
	.A(\addr_calc/fir_write_addr[25] ));
   TBUFX16TS \addr_calc/addr_tri6[31]  (.Y(addr[31]), 
	.OE(FE_OFN292_n2641), 
	.A(\addr_calc/iir_write_addr[31] ));
   TBUFX4TS \addr_calc/addr_tri3[17]  (.Y(addr[17]), 
	.OE(FE_OFN168_n195), 
	.A(\addr_calc/fir_read_addr[17] ));
   TBUFX4TS \addr_calc/addr_tri3[20]  (.Y(addr[20]), 
	.OE(FE_OFN169_n195), 
	.A(\addr_calc/fir_read_addr[20] ));
   TBUFX16TS \addr_calc/addr_tri2[25]  (.Y(addr[25]), 
	.OE(FE_OFN303_n2645), 
	.A(\addr_calc/fft_write_addr[25] ));
   TBUFX16TS \addr_calc/addr_tri6[25]  (.Y(addr[25]), 
	.OE(FE_OFN291_n2641), 
	.A(FE_OFN126_addr_calc_iir_write_addr_25_));
   TBUFX12TS \addr_calc/addr_tri6[28]  (.Y(addr[28]), 
	.OE(FE_OFN289_n2641), 
	.A(\addr_calc/iir_write_addr[28] ));
   TBUFX12TS \addr_calc/addr_tri3[27]  (.Y(addr[27]), 
	.OE(FE_OFN307_n2644), 
	.A(\addr_calc/fir_read_addr[27] ));
   TBUFX12TS \addr_calc/addr_tri[27]  (.Y(addr[27]), 
	.OE(FE_OFN299_n2646), 
	.A(\addr_calc/fft_read_addr[27] ));
   TBUFX12TS \addr_calc/addr_tri6[27]  (.Y(addr[27]), 
	.OE(FE_OFN291_n2641), 
	.A(\addr_calc/iir_write_addr[27] ));
   DFFHQX4TS \addr_calc/fir_read_calc/counter/count_reg[9]  (.Q(\addr_calc/fir_read_calc/count[9] ), 
	.D(n1089), 
	.CK(clk__L1_N0));
   TBUFX16TS \addr_calc/addr_tri2[23]  (.Y(addr[23]), 
	.OE(FE_OFN166_n259), 
	.A(\addr_calc/fft_write_addr[23] ));
   TBUFX16TS \addr_calc/addr_tri2[31]  (.Y(addr[31]), 
	.OE(FE_OFN304_n2645), 
	.A(\addr_calc/fft_write_addr[31] ));
   DFFHQX2TS \addr_calc/fft_read_calc/counter/count_reg[6]  (.Q(\addr_calc/fft_read_calc/count[6] ), 
	.D(n1028), 
	.CK(clk__L1_N0));
   TBUFX16TS \addr_calc/addr_tri2[27]  (.Y(addr[27]), 
	.OE(FE_OFN303_n2645), 
	.A(\addr_calc/fft_write_addr[27] ));
   TBUFX16TS \addr_calc/addr_tri5[29]  (.Y(addr[29]), 
	.OE(FE_OFN296_n2642), 
	.A(\addr_calc/iir_read_addr[29] ));
   NAND2X4TS U399 (.Y(\addr_calc/iir_write_calc/counter/N38 ), 
	.B(n1780), 
	.A(n1779));
   XNOR2X2TS U400 (.Y(\addr_calc/fir_write_addr[30] ), 
	.B(n1538), 
	.A(\add_x_19_3/n38 ));
   OAI21X2TS U401 (.Y(\add_x_19_4/n99 ), 
	.B0(\add_x_19_4/n101 ), 
	.A1(\add_x_19_4/n102 ), 
	.A0(\add_x_19_4/n100 ));
   XNOR2X1TS U402 (.Y(\DP_OP_158_296_6262/n202 ), 
	.B(n1988), 
	.A(\DP_OP_158_296_6262/n841 ));
   NOR2X4TS U404 (.Y(\add_x_19_0/n84 ), 
	.B(\add_x_19_0/n89 ), 
	.A(\add_x_19_0/n86 ));
   XOR2X4TS U405 (.Y(\addr_calc/fir_read_addr[19] ), 
	.B(n1137), 
	.A(\add_x_19_2/n99 ));
   AND2X4TS U406 (.Y(n1137), 
	.B(\add_x_19_2/n98 ), 
	.A(\add_x_19_2/n204 ));
   XOR2XLTS U407 (.Y(\DP_OP_159_297_3515/n495 ), 
	.B(n1971), 
	.A(n1702));
   NAND2X2TS U408 (.Y(\add_x_19_0/n90 ), 
	.B(n2441), 
	.A(\addr_calc/fft_read_calc/count[20] ));
   NOR2XLTS U409 (.Y(n1138), 
	.B(FE_OFN491_filesize_9_), 
	.A(FE_OFN492_filesize_8_));
   AO22X1TS U411 (.Y(n1105), 
	.B1(FE_OCPUNCON1088_n2805), 
	.B0(\addr_calc/fir_write_calc/count[25] ), 
	.A1(\addr_calc/fir_write_calc/counter/N68 ), 
	.A0(FE_OFN50_n2803));
   INVX12TS U413 (.Y(n1758), 
	.A(FE_OFN49_n2803));
   NOR2X1TS U414 (.Y(n2803), 
	.B(n785), 
	.A(n1241));
   INVX3TS U415 (.Y(\add_x_19_1/n91 ), 
	.A(\add_x_19_1/n92 ));
   XOR2X4TS U418 (.Y(\addr_calc/fft_write_addr[24] ), 
	.B(n1406), 
	.A(FE_OCP_RBN1379_add_x_19_1_n69));
   OAI21X2TS U419 (.Y(\add_x_19_1/n57 ), 
	.B0(\add_x_19_1/n59 ), 
	.A1(\add_x_19_1/n58 ), 
	.A0(\add_x_19_1/n60 ));
   OAI2BB1X2TS U421 (.Y(n1028), 
	.B0(n1608), 
	.A1N(FE_OFN14_n2794), 
	.A0N(\addr_calc/fft_read_calc/count[6] ));
   XOR2X4TS U424 (.Y(\addr_calc/fft_read_addr[20] ), 
	.B(n1393), 
	.A(FE_OCP_RBN1383_add_x_19_0_n92));
   MXI2X1TS U425 (.Y(n1066), 
	.S0(n2797), 
	.B(\addr_calc/fft_write_calc/counter/N43 ), 
	.A(n2798));
   XOR2X1TS U426 (.Y(\DP_OP_158_296_6262/n580 ), 
	.B(\add_x_22_1/n30 ), 
	.A(n1731));
   XOR2X4TS U427 (.Y(\addr_calc/fir_read_addr[26] ), 
	.B(n1325), 
	.A(\add_x_19_2/n60 ));
   XOR2XLTS U429 (.Y(\addr_calc/fir_read_addr[8] ), 
	.B(\add_x_19_2/n24 ), 
	.A(\add_x_19_2/n156 ));
   XOR2X4TS U430 (.Y(\addr_calc/fir_write_addr[31] ), 
	.B(n1140), 
	.A(\add_x_19_3/n35 ));
   AND2X6TS U431 (.Y(n1140), 
	.B(\add_x_19_3/n34 ), 
	.A(n2630));
   INVX2TS U432 (.Y(n1751), 
	.A(n1701));
   NAND2X1TS U433 (.Y(n1141), 
	.B(\addr_calc/fir_read_calc/counter/N47 ), 
	.A(FE_OFN61_n2807));
   NAND2X1TS U434 (.Y(n1142), 
	.B(n1906), 
	.A(FE_OFN71_n2809));
   NAND2X1TS U435 (.Y(n1094), 
	.B(n1142), 
	.A(n1141));
   NOR2X1TS U438 (.Y(\DP_OP_159_297_3515/n1011 ), 
	.B(\DP_OP_159_297_3515/n1014 ), 
	.A(\DP_OP_159_297_3515/n1026 ));
   CLKINVX2TS U440 (.Y(n1540), 
	.A(n1897));
   NAND4BX2TS U441 (.Y(\add_x_22_2/n94 ), 
	.D(n2001), 
	.C(FE_OFN227_addr_calc_fir_read_calc_count_7_), 
	.B(\add_x_22_2/n111 ), 
	.AN(\add_x_22_2/n103 ));
   XNOR2X4TS U442 (.Y(\addr_calc/fir_read_addr[23] ), 
	.B(n1597), 
	.A(n1596));
   OAI21X2TS U443 (.Y(\add_x_19_1/n80 ), 
	.B0(\add_x_19_1/n82 ), 
	.A1(\add_x_19_1/n81 ), 
	.A0(\add_x_19_1/n83 ));
   NOR4BBX1TS U444 (.Y(n877), 
	.D(n2001), 
	.C(FE_OFN227_addr_calc_fir_read_calc_count_7_), 
	.BN(n1143), 
	.AN(n1899));
   CLKINVX2TS U445 (.Y(n1143), 
	.A(n1997));
   AOI2BB1X2TS U446 (.Y(\addr_calc/fir_read_addr[27] ), 
	.B0(n1228), 
	.A1N(n1227), 
	.A0N(\add_x_19_2/n60 ));
   AOI21X4TS U447 (.Y(\add_x_19_1/n60 ), 
	.B0(\add_x_19_1/n62 ), 
	.A1(\add_x_19_1/n61 ), 
	.A0(\add_x_19_1/n69 ));
   NOR2X4TS U452 (.Y(\add_x_19_3/n86 ), 
	.B(FE_OCPUNCON1078_FE_OFN377_offset_21_), 
	.A(n1892));
   CLKINVX2TS U453 (.Y(n1892), 
	.A(n1891));
   AND2X2TS U454 (.Y(n1698), 
	.B(\DP_OP_159_297_3515/n963 ), 
	.A(n1789));
   CLKINVX2TS U455 (.Y(n2048), 
	.A(n2047));
   NOR2X2TS U456 (.Y(\DP_OP_159_297_3515/n956 ), 
	.B(\DP_OP_159_297_3515/n959 ), 
	.A(\DP_OP_159_297_3515/n971 ));
   XOR2X1TS U457 (.Y(n1659), 
	.B(\DP_OP_159_297_3515/n871 ), 
	.A(\DP_OP_158_296_6262/n1950 ));
   CLKINVX2TS U458 (.Y(\DP_OP_159_297_3515/n871 ), 
	.A(FE_OFN487_filesize_13_));
   XNOR2X1TS U459 (.Y(\DP_OP_159_297_3515/n289 ), 
	.B(FE_OFN248_addr_calc_iir_read_calc_count_10_), 
	.A(n2621));
   NOR2X1TS U460 (.Y(\DP_OP_159_297_3515/n1040 ), 
	.B(\DP_OP_159_297_3515/n1041 ), 
	.A(\DP_OP_159_297_3515/n1052 ));
   NAND2X1TS U461 (.Y(\DP_OP_158_296_6262/n318 ), 
	.B(\DP_OP_158_296_6262/n347 ), 
	.A(\DP_OP_158_296_6262/n320 ));
   NOR2X1TS U462 (.Y(\DP_OP_158_296_6262/n1158 ), 
	.B(\DP_OP_158_296_6262/n1160 ), 
	.A(\DP_OP_158_296_6262/n1171 ));
   CLKINVX6TS U463 (.Y(n1789), 
	.A(n1782));
   CLKINVX4TS U464 (.Y(\add_x_19_4/n91 ), 
	.A(\add_x_19_4/n92 ));
   XNOR2XLTS U467 (.Y(n1634), 
	.B(\addr_calc/fft_read_calc/count[17] ), 
	.A(n1635));
   INVXLTS U468 (.Y(\add_x_19_0/n206 ), 
	.A(\add_x_19_0/n105 ));
   XNOR2X2TS U469 (.Y(\DP_OP_159_297_3515/n5 ), 
	.B(FE_OFN234_addr_calc_iir_read_calc_count_31_), 
	.A(n2614));
   XOR2X4TS U470 (.Y(n1738), 
	.B(n1146), 
	.A(\DP_OP_159_297_3515/n934 ));
   CLKINVX2TS U471 (.Y(n1146), 
	.A(\DP_OP_158_296_6262/n1869 ));
   XNOR2X1TS U472 (.Y(\DP_OP_158_296_6262/n724 ), 
	.B(n2023), 
	.A(n1756));
   AOI21X2TS U473 (.Y(\add_x_19_1/n167 ), 
	.B0(n1157), 
	.A1(\add_x_19_1/n168 ), 
	.A0(\add_x_19_1/n177 ));
   NOR2X4TS U474 (.Y(\add_x_19_3/n131 ), 
	.B(FE_OFN232_addr_calc_fir_write_calc_count_12_), 
	.A(FE_OFN413_offset_12_));
   OAI21X4TS U476 (.Y(\add_x_19_3/n65 ), 
	.B0(\add_x_19_3/n67 ), 
	.A1(\add_x_19_3/n66 ), 
	.A0(\add_x_19_3/n68 ));
   XNOR2X4TS U479 (.Y(\addr_calc/iir_read_addr[31] ), 
	.B(n1357), 
	.A(n1356));
   NAND2XLTS U480 (.Y(\DP_OP_158_296_6262/n1944 ), 
	.B(\DP_OP_158_296_6262/n1945 ), 
	.A(\DP_OP_158_296_6262/n1959 ));
   OAI21XLTS U481 (.Y(n1394), 
	.B0(fft_enable), 
	.A1(n2057), 
	.A0(n2793));
   NOR2BX4TS U483 (.Y(\add_x_19_4/n126 ), 
	.B(\add_x_19_4/n131 ), 
	.AN(n1632));
   OAI21X2TS U485 (.Y(\add_x_19_4/n127 ), 
	.B0(\add_x_19_4/n129 ), 
	.A1(\add_x_19_4/n128 ), 
	.A0(\add_x_19_4/n132 ));
   XNOR2X1TS U486 (.Y(\DP_OP_158_296_6262/n621 ), 
	.B(FE_OFN281_addr_calc_fft_write_calc_count_20_), 
	.A(n1776));
   NAND2X1TS U487 (.Y(n1147), 
	.B(n1462), 
	.A(n1677));
   CLKINVX2TS U491 (.Y(\DP_OP_158_296_6262/n1959 ), 
	.A(\DP_OP_158_296_6262/n1958 ));
   XOR2X1TS U492 (.Y(\DP_OP_158_296_6262/n39 ), 
	.B(n1841), 
	.A(n1463));
   OAI21X1TS U493 (.Y(\add_x_19_3/n50 ), 
	.B0(\add_x_19_3/n52 ), 
	.A1(\add_x_19_3/n51 ), 
	.A0(\add_x_19_3/n68 ));
   NAND2X4TS U495 (.Y(\DP_OP_158_296_6262/n1958 ), 
	.B(n1591), 
	.A(\DP_OP_158_296_6262/n1973 ));
   XOR2X4TS U496 (.Y(\addr_calc/fft_read_addr[27] ), 
	.B(n1465), 
	.A(\add_x_19_0/n57 ));
   XNOR2X1TS U497 (.Y(\DP_OP_158_296_6262/n1136 ), 
	.B(\addr_calc/fft_read_calc/count[15] ), 
	.A(n1658));
   NOR2X1TS U498 (.Y(\DP_OP_158_296_6262/n996 ), 
	.B(\DP_OP_158_296_6262/n1013 ), 
	.A(\DP_OP_158_296_6262/n998 ));
   MXI2X4TS U499 (.Y(\DP_OP_159_297_3515/n1064 ), 
	.S0(\DP_OP_159_297_3515/n1075 ), 
	.B(\DP_OP_159_297_3515/n1066 ), 
	.A(\DP_OP_159_297_3515/n880 ));
   XNOR2X1TS U500 (.Y(\DP_OP_159_297_3515/n705 ), 
	.B(n1942), 
	.A(n2620));
   NAND2X1TS U501 (.Y(n2620), 
	.B(n1735), 
	.A(n1734));
   NOR2X4TS U502 (.Y(\DP_OP_158_296_6262/n1878 ), 
	.B(FE_OFN473_filesize_23_), 
	.A(FE_OFN475_filesize_22_));
   NOR2X1TS U504 (.Y(\DP_OP_158_296_6262/n687 ), 
	.B(\DP_OP_158_296_6262/n689 ), 
	.A(\DP_OP_158_296_6262/n702 ));
   XNOR2X1TS U506 (.Y(\DP_OP_158_296_6262/n1216 ), 
	.B(n1666), 
	.A(n1651));
   NOR2X2TS U507 (.Y(\add_x_19_4/n123 ), 
	.B(\addr_calc/iir_read_calc/count[14] ), 
	.A(FE_OFN405_offset_14_));
   NOR2X2TS U508 (.Y(\add_x_19_4/n139 ), 
	.B(FE_OFN417_offset_11_), 
	.A(FE_OFN237_addr_calc_iir_read_calc_count_11_));
   CLKXOR2X8TS U509 (.Y(n1655), 
	.B(FE_OFN470_filesize_25_), 
	.A(n1147));
   NOR2X8TS U510 (.Y(\DP_OP_158_296_6262/n1945 ), 
	.B(FE_OFN488_filesize_12_), 
	.A(FE_OFN487_filesize_13_));
   OAI31X4TS U511 (.Y(\addr_calc/fir_write_addr[13] ), 
	.B0(n1302), 
	.A2(n1301), 
	.A1(n1300), 
	.A0(\add_x_19_3/n128 ));
   XNOR2X4TS U513 (.Y(\addr_calc/iir_read_addr[28] ), 
	.B(\add_x_19_4/n4 ), 
	.A(\add_x_19_4/n50 ));
   XNOR2X4TS U514 (.Y(\addr_calc/iir_read_addr[25] ), 
	.B(\add_x_19_4/n7 ), 
	.A(\add_x_19_4/n65 ));
   NAND4X2TS U515 (.Y(n2799), 
	.D(n879), 
	.C(n878), 
	.B(n877), 
	.A(n876));
   NOR4X1TS U516 (.Y(n879), 
	.D(n1871), 
	.C(n1842), 
	.B(n2004), 
	.A(n1838));
   CLKINVX2TS U517 (.Y(n1871), 
	.A(n1870));
   NOR2X8TS U518 (.Y(\add_x_19_5/n162 ), 
	.B(n1683), 
	.A(FE_OCP_RBN1840_offset_7_));
   INVX4TS U519 (.Y(n1683), 
	.A(n1938));
   OAI21X2TS U520 (.Y(\add_x_19_0/n57 ), 
	.B0(\add_x_19_0/n59 ), 
	.A1(\add_x_19_0/n58 ), 
	.A0(\add_x_19_0/n60 ));
   NOR2X2TS U521 (.Y(\DP_OP_158_296_6262/n513 ), 
	.B(\DP_OP_158_296_6262/n534 ), 
	.A(\DP_OP_158_296_6262/n515 ));
   NAND2X2TS U522 (.Y(\add_x_19_1/n171 ), 
	.B(FE_OCP_RBN1494_offset_5_), 
	.A(\addr_calc/fft_write_calc/count[5] ));
   XOR2X1TS U523 (.Y(\addr_calc/fft_write_addr[8] ), 
	.B(n1405), 
	.A(FE_OCP_RBN1956_FE_OFN520_add_x_19_1_n157));
   XNOR2X4TS U525 (.Y(\addr_calc/fft_write_addr[10] ), 
	.B(\add_x_19_1/n146 ), 
	.A(n1446));
   NOR2X2TS U526 (.Y(\add_x_19_3/n97 ), 
	.B(FE_OCPUNCON1079_FE_OFN382_offset_19_), 
	.A(n1670));
   CLKINVX2TS U527 (.Y(n1670), 
	.A(n1889));
   NOR2X8TS U528 (.Y(\add_x_19_5/n170 ), 
	.B(n1686), 
	.A(FE_OCP_RBN1492_offset_5_));
   XNOR2X4TS U529 (.Y(\addr_calc/fir_write_addr[23] ), 
	.B(\add_x_19_3/n9 ), 
	.A(\add_x_19_3/n80 ));
   NAND2XLTS U530 (.Y(\add_x_22_3/n65 ), 
	.B(\addr_calc/fir_write_calc/count[14] ), 
	.A(\add_x_22_3/n68 ));
   NAND4BXLTS U532 (.Y(n1273), 
	.D(\add_x_22_3/n77 ), 
	.C(n1883), 
	.B(n2003), 
	.AN(\add_x_22_3/n69 ));
   CLKINVX2TS U534 (.Y(n2002), 
	.A(\addr_calc/fir_write_calc/count[14] ));
   CLKINVX2TS U536 (.Y(n1889), 
	.A(\addr_calc/fir_write_calc/count[19] ));
   CLKINVX2TS U537 (.Y(\add_x_22_0/n40 ), 
	.A(\addr_calc/fft_read_calc/count[20] ));
   NOR2BX2TS U538 (.Y(\add_x_19_0/n89 ), 
	.B(\addr_calc/fft_read_calc/count[20] ), 
	.AN(FE_OCP_RBN1363_FE_OCP_DRV_N1167_offset_20_));
   NOR2X6TS U539 (.Y(\add_x_19_4/n162 ), 
	.B(FE_OFN247_addr_calc_iir_read_calc_count_7_), 
	.A(FE_OCP_RBN1840_offset_7_));
   CLKINVX2TS U540 (.Y(n1158), 
	.A(\addr_calc/fft_write_calc/count[5] ));
   NOR2X2TS U541 (.Y(\DP_OP_158_296_6262/n1978 ), 
	.B(n2364), 
	.A(n1728));
   NOR2X2TS U542 (.Y(\DP_OP_158_296_6262/n1971 ), 
	.B(\DP_OP_158_296_6262/n1972 ), 
	.A(n1728));
   NOR2X2TS U543 (.Y(\DP_OP_158_296_6262/n1936 ), 
	.B(\DP_OP_158_296_6262/n1937 ), 
	.A(n1728));
   CLKINVX2TS U544 (.Y(\DP_OP_159_297_3515/n875 ), 
	.A(FE_OFN491_filesize_9_));
   CLKINVX2TS U547 (.Y(n1900), 
	.A(n1899));
   XOR2X4TS U549 (.Y(n1149), 
	.B(n1678), 
	.A(FE_OCPN1910_n1736));
   XOR2X1TS U551 (.Y(\DP_OP_158_296_6262/n534 ), 
	.B(\add_x_22_1/n15 ), 
	.A(\DP_OP_158_296_6262/n833 ));
   XNOR2X2TS U552 (.Y(\addr_calc/fft_write_addr[26] ), 
	.B(n1150), 
	.A(\add_x_19_1/n60 ));
   CLKINVX2TS U553 (.Y(n1150), 
	.A(n1321));
   AO22X1TS U555 (.Y(n1082), 
	.B1(\addr_calc/fir_read_calc/count[16] ), 
	.B0(FE_OFN64_n2809), 
	.A1(\addr_calc/fir_read_calc/counter/N59 ), 
	.A0(FE_OFN53_n2807));
   AO22X1TS U556 (.Y(n1080), 
	.B1(\addr_calc/fir_read_calc/count[18] ), 
	.B0(FE_OFN65_n2809), 
	.A1(\addr_calc/fir_read_calc/counter/N61 ), 
	.A0(FE_OFN55_n2807));
   NAND2BX2TS U557 (.Y(\add_x_19_5/n90 ), 
	.B(FE_OFN558_n2441), 
	.AN(n2047));
   NAND2XLTS U558 (.Y(\DP_OP_159_297_3515/n1041 ), 
	.B(FE_OFN492_filesize_8_), 
	.A(FE_OFN493_filesize_7_));
   XNOR2X1TS U559 (.Y(\DP_OP_159_297_3515/n269 ), 
	.B(n1785), 
	.A(n2619));
   OAI2BB1XLTS U563 (.Y(n1068), 
	.B0(n1645), 
	.A1N(\addr_calc/fir_read_calc/counter/N73 ), 
	.A0N(FE_OFN59_n2807));
   NAND2BXLTS U565 (.Y(n1188), 
	.B(FE_OFN60_n2807), 
	.AN(n1189));
   AO22X2TS U566 (.Y(n1091), 
	.B1(FE_OFN227_addr_calc_fir_read_calc_count_7_), 
	.B0(FE_OFN71_n2809), 
	.A1(\addr_calc/fir_read_calc/counter/N50 ), 
	.A0(FE_OFN61_n2807));
   NAND2BXLTS U567 (.Y(n1202), 
	.B(FE_OFN58_n2807), 
	.AN(n1203));
   AO22X1TS U568 (.Y(n1097), 
	.B1(\addr_calc/fir_read_calc/count[1] ), 
	.B0(FE_OFN66_n2809), 
	.A1(\addr_calc/fir_read_calc/counter/N44 ), 
	.A0(FE_OFN56_n2807));
   NAND2BX1TS U569 (.Y(n1167), 
	.B(FE_OFN58_n2807), 
	.AN(n1168));
   AO22X2TS U570 (.Y(n1093), 
	.B1(\addr_calc/fir_read_calc/count[5] ), 
	.B0(FE_OFN71_n2809), 
	.A1(\addr_calc/fir_read_calc/counter/N48 ), 
	.A0(FE_OFN61_n2807));
   NAND2BXLTS U571 (.Y(n1184), 
	.B(FE_OFN60_n2807), 
	.AN(n1185));
   INVX2TS U575 (.Y(n1754), 
	.A(n1701));
   OAI2BB1XLTS U578 (.Y(n1071), 
	.B0(n1202), 
	.A1N(FE_OFN68_n2809), 
	.A0N(\addr_calc/fir_read_calc/count[27] ));
   INVX8TS U579 (.Y(n1762), 
	.A(FE_OFN47_n1758));
   XNOR2X1TS U584 (.Y(\DP_OP_158_296_6262/n1042 ), 
	.B(n1665), 
	.A(n1652));
   NOR2X6TS U585 (.Y(\DP_OP_158_296_6262/n1906 ), 
	.B(FE_OFN478_filesize_19_), 
	.A(FE_OFN479_filesize_18_));
   NAND2X2TS U587 (.Y(\DP_OP_158_296_6262/n576 ), 
	.B(\DP_OP_158_296_6262/n578 ), 
	.A(\DP_OP_158_296_6262/n606 ));
   INVX1TS U588 (.Y(n1479), 
	.A(n1158));
   OAI21XLTS U589 (.Y(n1157), 
	.B0(\add_x_19_1/n171 ), 
	.A1(\add_x_19_1/n176 ), 
	.A0(\add_x_19_1/n170 ));
   AOI21X4TS U591 (.Y(\add_x_19_1/n113 ), 
	.B0(\add_x_19_1/n115 ), 
	.A1(\add_x_19_1/n114 ), 
	.A0(FE_OFN520_add_x_19_1_n157));
   OAI21X4TS U592 (.Y(\add_x_19_1/n92 ), 
	.B0(\add_x_19_1/n94 ), 
	.A1(\add_x_19_1/n93 ), 
	.A0(FE_OFN523_add_x_19_1_n113));
   INVX12TS U594 (.Y(\add_x_19_1/n112 ), 
	.A(FE_OFN523_add_x_19_1_n113));
   OAI21X4TS U595 (.Y(\add_x_19_1/n69 ), 
	.B0(\add_x_19_1/n71 ), 
	.A1(\add_x_19_1/n70 ), 
	.A0(FE_OFN523_add_x_19_1_n113));
   AOI21X4TS U596 (.Y(\add_x_19_1/n83 ), 
	.B0(\add_x_19_1/n85 ), 
	.A1(\add_x_19_1/n84 ), 
	.A0(\add_x_19_1/n92 ));
   XNOR2X2TS U597 (.Y(\addr_calc/fft_write_addr[22] ), 
	.B(n1154), 
	.A(\add_x_19_1/n83 ));
   NAND2BX1TS U598 (.Y(n1153), 
	.B(\add_x_19_1/n82 ), 
	.AN(\add_x_19_1/n81 ));
   INVX2TS U599 (.Y(n1154), 
	.A(n1153));
   NAND2X1TS U600 (.Y(\DP_OP_158_296_6262/n1998 ), 
	.B(\DP_OP_158_296_6262/n1999 ), 
	.A(\DP_OP_158_296_6262/n2010 ));
   INVX2TS U601 (.Y(n1155), 
	.A(FE_OFN469_filesize_25_));
   NOR2X4TS U602 (.Y(\add_x_19_4/n120 ), 
	.B(FE_OCPUNCON1942_FE_OFN399_offset_15_), 
	.A(\addr_calc/iir_read_calc/count[15] ));
   INVXLTS U603 (.Y(\add_x_19_1/n218 ), 
	.A(\add_x_19_1/n170 ));
   XNOR2X4TS U604 (.Y(\addr_calc/iir_read_addr[22] ), 
	.B(n1156), 
	.A(\add_x_19_4/n83 ));
   CLKINVX2TS U605 (.Y(n1156), 
	.A(n1433));
   XOR2X1TS U607 (.Y(n1602), 
	.B(FE_OFN251_addr_calc_fft_read_calc_count_5_), 
	.A(n2595));
   XNOR2X1TS U608 (.Y(\DP_OP_159_297_3515/n638 ), 
	.B(n1954), 
	.A(n2607));
   OR3X1TS U609 (.Y(n1737), 
	.C(n1860), 
	.B(n2785), 
	.A(FE_OFN326_data_cntl_N191));
   NOR2X8TS U610 (.Y(n1781), 
	.B(\DP_OP_159_297_3515/n160 ), 
	.A(\DP_OP_159_297_3515/n1 ));
   XOR2XLTS U612 (.Y(\DP_OP_159_297_3515/n625 ), 
	.B(FE_OFN266_addr_calc_iir_write_calc_count_18_), 
	.A(\DP_OP_159_297_3515/n1128 ));
   NOR2X4TS U613 (.Y(\DP_OP_158_296_6262/n1933 ), 
	.B(FE_OFN486_filesize_14_), 
	.A(FE_OFN484_filesize_15_));
   XNOR2X4TS U615 (.Y(\addr_calc/iir_write_addr[28] ), 
	.B(\add_x_19_5/n4 ), 
	.A(\add_x_19_5/n50 ));
   NAND2BX1TS U616 (.Y(\add_x_22_1/n103 ), 
	.B(n1939), 
	.AN(n1158));
   AOI21X4TS U617 (.Y(\add_x_19_1/n159 ), 
	.B0(\add_x_19_1/n161 ), 
	.A1(\add_x_19_1/n160 ), 
	.A0(\add_x_19_1/n169 ));
   NAND2X2TS U620 (.Y(\add_x_19_1/n158 ), 
	.B(\add_x_19_1/n168 ), 
	.A(\add_x_19_1/n160 ));
   XNOR2X1TS U621 (.Y(n1159), 
	.B(n1912), 
	.A(n1161));
   NOR2BX1TS U622 (.Y(n1161), 
	.B(n1162), 
	.AN(\add_x_22_1/n16 ));
   CLKINVX2TS U623 (.Y(n1162), 
	.A(n2574));
   NAND2X1TS U624 (.Y(n1160), 
	.B(\addr_calc/fft_write_calc/count[27] ), 
	.A(FE_OFN23_n2797));
   OAI2BB1X1TS U625 (.Y(n1039), 
	.B0(n1160), 
	.A1N(n1159), 
	.A0N(FE_OFN32_n2795));
   XNOR2X1TS U626 (.Y(n1164), 
	.B(FE_OFN276_addr_calc_fft_write_calc_count_24_), 
	.A(\add_x_22_1/n23 ));
   NAND2BX1TS U628 (.Y(n1163), 
	.B(FE_OFN31_n2795), 
	.AN(n1164));
   OAI2BB1X1TS U629 (.Y(n1042), 
	.B0(n1163), 
	.A1N(\addr_calc/fft_write_calc/count[24] ), 
	.A0N(FE_OFN22_n2797));
   NAND2X1TS U630 (.Y(n1166), 
	.B(\addr_calc/fft_write_calc/counter/N69 ), 
	.A(FE_OFN32_n2795));
   OAI2BB1X1TS U631 (.Y(n1040), 
	.B0(n1166), 
	.A1N(FE_OFN23_n2797), 
	.A0N(n2574));
   XNOR2X1TS U632 (.Y(n1168), 
	.B(n1875), 
	.A(n1169));
   NAND2BX1TS U633 (.Y(n1169), 
	.B(\add_x_22_2/n23 ), 
	.AN(n1170));
   CLKINVX2TS U634 (.Y(n1170), 
	.A(\addr_calc/fir_read_calc/count[24] ));
   OAI2BB1X1TS U635 (.Y(n1073), 
	.B0(n1167), 
	.A1N(FE_OFN68_n2809), 
	.A0N(\addr_calc/fir_read_calc/count[25] ));
   XNOR2X1TS U636 (.Y(n1172), 
	.B(\addr_calc/fir_write_calc/count[26] ), 
	.A(\add_x_22_3/n16 ));
   NAND2BX1TS U638 (.Y(n1171), 
	.B(FE_OFN549_n1763), 
	.AN(n1172));
   OAI2BB1X1TS U639 (.Y(n1104), 
	.B0(n1171), 
	.A1N(FE_OCPUNCON1089_n2805), 
	.A0N(\addr_calc/fir_write_calc/count[26] ));
   CLKINVX1TS U640 (.Y(\add_x_19_1/n204 ), 
	.A(\add_x_19_1/n97 ));
   OAI21X1TS U641 (.Y(\add_x_19_1/n99 ), 
	.B0(\add_x_19_1/n101 ), 
	.A1(\add_x_19_1/n100 ), 
	.A0(\add_x_19_1/n102 ));
   XNOR2X2TS U642 (.Y(\addr_calc/fft_write_addr[19] ), 
	.B(\add_x_19_1/n13 ), 
	.A(\add_x_19_1/n99 ));
   OAI2BB1X1TS U643 (.Y(n1177), 
	.B0(n1179), 
	.A1N(n1178), 
	.A0N(FE_OFN143_add_x_19_3_n59));
   OAI2BB1X1TS U644 (.Y(n1179), 
	.B0(n1180), 
	.A1N(FE_OFN143_add_x_19_3_n59), 
	.A0N(\add_x_19_3/n58 ));
   CLKINVX2TS U645 (.Y(n1180), 
	.A(n1178));
   NOR2BX1TS U646 (.Y(n1176), 
	.B(n1178), 
	.AN(FE_OFN143_add_x_19_3_n59));
   NAND2BX1TS U647 (.Y(n1174), 
	.B(n1178), 
	.AN(\add_x_19_3/n58 ));
   NOR2BX1TS U648 (.Y(n1178), 
	.B(\add_x_19_3/n55 ), 
	.AN(\add_x_19_3/n56 ));
   AOI2BB1X4TS U649 (.Y(\addr_calc/fir_write_addr[27] ), 
	.B0(n1175), 
	.A1N(n1174), 
	.A0N(\add_x_19_3/n60 ));
   OAI2BB1X2TS U650 (.Y(n1175), 
	.B0(n1177), 
	.A1N(\add_x_19_3/n60 ), 
	.A0N(n1176));
   XNOR2X1TS U651 (.Y(n1182), 
	.B(\addr_calc/iir_write_calc/count[18] ), 
	.A(\add_x_22_5/n50 ));
   NAND2BX1TS U653 (.Y(n1181), 
	.B(FE_OCPUNCON1882_n2813), 
	.AN(n1182));
   OAI2BB1X1TS U654 (.Y(n984), 
	.B0(n1181), 
	.A1N(FE_OCPUNCON1571_n2812), 
	.A0N(\addr_calc/iir_write_calc/count[18] ));
   AO22X1TS U655 (.Y(n982), 
	.B1(\addr_calc/iir_write_calc/count[20] ), 
	.B0(FE_OCPUNCON1571_n2812), 
	.A1(\addr_calc/iir_write_calc/counter/N63 ), 
	.A0(FE_OCPUNCON1883_n2813));
   XNOR2X1TS U656 (.Y(n1185), 
	.B(\add_x_22_2/n114 ), 
	.A(n1186));
   NAND2BX1TS U657 (.Y(n1186), 
	.B(\add_x_22_2/n118 ), 
	.AN(n1187));
   CLKINVX2TS U658 (.Y(n1187), 
	.A(n2004));
   OAI2BB1X1TS U659 (.Y(n1095), 
	.B0(n1184), 
	.A1N(FE_OFN70_n2809), 
	.A0N(n1908));
   AO22X1TS U660 (.Y(n1083), 
	.B1(n1890), 
	.B0(FE_OFN64_n2809), 
	.A1(\addr_calc/fir_read_calc/counter/N58 ), 
	.A0(FE_OFN53_n2807));
   XNOR2X1TS U661 (.Y(n1189), 
	.B(\addr_calc/fir_read_calc/count[31] ), 
	.A(\add_x_22_2/n1 ));
   OAI2BB1XLTS U662 (.Y(n1132), 
	.B0(n1188), 
	.A1N(FE_OFN70_n2809), 
	.A0N(\addr_calc/fir_read_calc/count[31] ));
   CLKINVX2TS U663 (.Y(n1191), 
	.A(\addr_calc/fir_write_calc/counter/N58 ));
   NAND2BX1TS U664 (.Y(n1190), 
	.B(FE_OFN548_n1763), 
	.AN(n1191));
   OAI2BB1X1TS U665 (.Y(n1115), 
	.B0(n1190), 
	.A1N(FE_OCPUNCON1085_n2805), 
	.A0N(\addr_calc/fir_write_calc/count[15] ));
   NOR2X4TS U666 (.Y(\add_x_19_2/n160 ), 
	.B(\add_x_19_2/n165 ), 
	.A(\add_x_19_2/n162 ));
   OAI21X2TS U667 (.Y(\add_x_19_2/n115 ), 
	.B0(\add_x_19_2/n117 ), 
	.A1(\add_x_19_2/n116 ), 
	.A0(\add_x_19_2/n136 ));
   AOI21X4TS U668 (.Y(\add_x_19_2/n113 ), 
	.B0(\add_x_19_2/n115 ), 
	.A1(\add_x_19_2/n114 ), 
	.A0(FE_OFN122_add_x_19_2_n157));
   INVX2TS U669 (.Y(\add_x_19_2/n71 ), 
	.A(\add_x_19_2/n73 ));
   INVX2TS U670 (.Y(\add_x_19_2/n70 ), 
	.A(\add_x_19_2/n72 ));
   OAI21X4TS U671 (.Y(\add_x_19_2/n69 ), 
	.B0(\add_x_19_2/n71 ), 
	.A1(\add_x_19_2/n70 ), 
	.A0(FE_OFN526_add_x_19_2_n113));
   CLKINVX1TS U672 (.Y(\add_x_19_2/n198 ), 
	.A(\add_x_19_2/n63 ));
   XNOR2X4TS U673 (.Y(\addr_calc/fir_read_addr[25] ), 
	.B(\add_x_19_2/n7 ), 
	.A(\add_x_19_2/n65 ));
   INVX1TS U674 (.Y(\add_x_19_2/n195 ), 
	.A(\add_x_19_2/n48 ));
   XNOR2X2TS U675 (.Y(\addr_calc/fir_read_addr[28] ), 
	.B(\add_x_19_2/n4 ), 
	.A(\add_x_19_2/n50 ));
   AOI21X1TS U676 (.Y(n2654), 
	.B0(n1860), 
	.A1(FE_OFN327_data_to_iir), 
	.A0(\addr_calc/iir_read_calc/counter/N38 ));
   AOI21X1TS U677 (.Y(n1192), 
	.B0(n1860), 
	.A1(FE_OFN327_data_to_iir), 
	.A0(\addr_calc/iir_read_calc/counter/N38 ));
   AO22X2TS U682 (.Y(n965), 
	.B1(n2018), 
	.B0(FE_OFN93_n1192), 
	.A1(\addr_calc/iir_read_calc/counter/N49 ), 
	.A0(FE_OFN84_n2787));
   AO22X1TS U683 (.Y(n967), 
	.B1(\addr_calc/iir_read_calc/count[4] ), 
	.B0(FE_OFN93_n1192), 
	.A1(\addr_calc/iir_read_calc/counter/N47 ), 
	.A0(FE_OFN84_n2787));
   AO22X1TS U684 (.Y(n968), 
	.B1(\addr_calc/iir_read_calc/count[3] ), 
	.B0(FE_OFN92_n1192), 
	.A1(\addr_calc/iir_read_calc/counter/N46 ), 
	.A0(FE_OFN83_n2787));
   AO22X2TS U685 (.Y(n966), 
	.B1(n2553), 
	.B0(FE_OFN93_n1192), 
	.A1(\addr_calc/iir_read_calc/counter/N48 ), 
	.A0(FE_OFN84_n2787));
   CLKINVX2TS U686 (.Y(n1195), 
	.A(\addr_calc/iir_read_calc/counter/N64 ));
   NAND2BX1TS U687 (.Y(n1194), 
	.B(FE_OFN79_n2787), 
	.AN(n1195));
   OAI2BB1X1TS U688 (.Y(n950), 
	.B0(n1194), 
	.A1N(FE_OFN87_n2654), 
	.A0N(\addr_calc/iir_read_calc/count[21] ));
   NAND2BX1TS U689 (.Y(n1196), 
	.B(FE_OFN86_n2654), 
	.AN(n2786));
   OAI21X1TS U690 (.Y(n971), 
	.B0(n1196), 
	.A1(FE_OFN86_n2654), 
	.A0(n1250));
   NAND2X4TS U691 (.Y(\DP_OP_159_297_3515/n1014 ), 
	.B(FE_OFN488_filesize_12_), 
	.A(FE_OFN489_filesize_11_));
   XNOR2X1TS U692 (.Y(n1198), 
	.B(n1200), 
	.A(n1199));
   CLKINVX2TS U693 (.Y(n1200), 
	.A(\add_x_22_4/n30 ));
   NOR2BX1TS U694 (.Y(n1199), 
	.B(n1201), 
	.AN(\add_x_22_4/n34 ));
   CLKINVX2TS U695 (.Y(n1201), 
	.A(n2031));
   NAND2BX1TS U696 (.Y(n1197), 
	.B(FE_OFN80_n2787), 
	.AN(n1198));
   OAI2BB1X1TS U697 (.Y(n948), 
	.B0(n1197), 
	.A1N(FE_OFN87_n2654), 
	.A0N(n2565));
   XNOR2X1TS U698 (.Y(n1203), 
	.B(FE_OFN243_addr_calc_fir_read_calc_count_27_), 
	.A(n1204));
   NOR2BX1TS U700 (.Y(n1204), 
	.B(n1206), 
	.AN(\add_x_22_2/n16 ));
   CLKINVX2TS U701 (.Y(n1206), 
	.A(FE_OFN270_addr_calc_fir_read_calc_count_26_));
   NAND2X1TS U702 (.Y(n1207), 
	.B(\addr_calc/fft_write_calc/counter/N61 ), 
	.A(FE_OFN29_n2795));
   OAI2BB1X1TS U703 (.Y(n1048), 
	.B0(n1207), 
	.A1N(FE_OFN20_n2797), 
	.A0N(\addr_calc/fft_write_calc/count[18] ));
   NOR2X1TS U704 (.Y(\DP_OP_158_296_6262/n1888 ), 
	.B(\DP_OP_158_296_6262/n1889 ), 
	.A(FE_OCPUNCON1081_n2589));
   XNOR2X4TS U705 (.Y(n1652), 
	.B(FE_OFN475_filesize_22_), 
	.A(\DP_OP_158_296_6262/n1888 ));
   XNOR2X1TS U706 (.Y(\DP_OP_158_296_6262/n822 ), 
	.B(\addr_calc/fft_write_calc/count[0] ), 
	.A(FE_OFN518_n2372));
   XOR2X1TS U707 (.Y(n1208), 
	.B(n2032), 
	.A(n2596));
   XOR2X1TS U708 (.Y(n1211), 
	.B(\addr_calc/fft_write_calc/count[4] ), 
	.A(\DP_OP_158_296_6262/n855 ));
   XOR2X1TS U709 (.Y(n1210), 
	.B(n2568), 
	.A(FE_OFN75_n2599));
   XOR2X1TS U710 (.Y(n1209), 
	.B(FE_OFN272_addr_calc_fft_write_calc_count_6_), 
	.A(n2593));
   XOR2X1TS U711 (.Y(n1212), 
	.B(n1479), 
	.A(n2595));
   XOR2X1TS U712 (.Y(\DP_OP_158_296_6262/n486 ), 
	.B(n1852), 
	.A(n1463));
   XNOR2X1TS U713 (.Y(\DP_OP_158_296_6262/n566 ), 
	.B(FE_OFN276_addr_calc_fft_write_calc_count_24_), 
	.A(FE_OCPN1732_n1718));
   XOR2XLTS U714 (.Y(n1213), 
	.B(n1915), 
	.A(n1655));
   XNOR2X1TS U715 (.Y(\DP_OP_158_296_6262/n515 ), 
	.B(n1913), 
	.A(n2602));
   XNOR2X1TS U716 (.Y(\DP_OP_158_296_6262/n595 ), 
	.B(FE_OFN284_addr_calc_fft_write_calc_count_22_), 
	.A(n1652));
   XNOR2X1TS U717 (.Y(\DP_OP_158_296_6262/n608 ), 
	.B(n1918), 
	.A(FE_OFN529_DP_OP_158_296_6262_n838));
   XNOR2X1TS U718 (.Y(\DP_OP_158_296_6262/n733 ), 
	.B(n1667), 
	.A(n1660));
   XNOR2X1TS U719 (.Y(\DP_OP_158_296_6262/n689 ), 
	.B(n1658), 
	.A(n1976));
   XNOR2X1TS U720 (.Y(\DP_OP_158_296_6262/n702 ), 
	.B(\addr_calc/fft_write_calc/count[14] ), 
	.A(n1657));
   XNOR2X1TS U721 (.Y(\DP_OP_158_296_6262/n664 ), 
	.B(\addr_calc/fft_write_calc/count[17] ), 
	.A(n1729));
   XOR2X1TS U722 (.Y(\DP_OP_158_296_6262/n649 ), 
	.B(n2019), 
	.A(\DP_OP_158_296_6262/n841 ));
   XNOR2X1TS U723 (.Y(\DP_OP_158_296_6262/n632 ), 
	.B(n1922), 
	.A(n1654));
   XOR2X1TS U724 (.Y(n1216), 
	.B(FE_OFN279_addr_calc_fft_write_calc_count_30_), 
	.A(\DP_OP_158_296_6262/n829 ));
   NOR2X1TS U725 (.Y(\DP_OP_158_296_6262/n484 ), 
	.B(\DP_OP_158_296_6262/n486 ), 
	.A(\DP_OP_158_296_6262/n501 ));
   NOR2BX1TS U726 (.Y(\DP_OP_158_296_6262/n549 ), 
	.B(\DP_OP_158_296_6262/n566 ), 
	.AN(n1213));
   NOR2X2TS U727 (.Y(\DP_OP_158_296_6262/n578 ), 
	.B(\DP_OP_158_296_6262/n580 ), 
	.A(\DP_OP_158_296_6262/n595 ));
   NOR2X2TS U728 (.Y(\DP_OP_158_296_6262/n606 ), 
	.B(\DP_OP_158_296_6262/n608 ), 
	.A(\DP_OP_158_296_6262/n621 ));
   NOR2X1TS U729 (.Y(\DP_OP_158_296_6262/n767 ), 
	.B(\DP_OP_158_296_6262/n776 ), 
	.A(\DP_OP_158_296_6262/n769 ));
   NOR2X1TS U730 (.Y(\DP_OP_158_296_6262/n751 ), 
	.B(\DP_OP_158_296_6262/n762 ), 
	.A(\DP_OP_158_296_6262/n753 ));
   NOR2X1TS U731 (.Y(\DP_OP_158_296_6262/n731 ), 
	.B(\DP_OP_158_296_6262/n733 ), 
	.A(\DP_OP_158_296_6262/n744 ));
   NOR2X1TS U732 (.Y(\DP_OP_158_296_6262/n711 ), 
	.B(\DP_OP_158_296_6262/n713 ), 
	.A(\DP_OP_158_296_6262/n724 ));
   NOR2X2TS U733 (.Y(\DP_OP_158_296_6262/n662 ), 
	.B(\DP_OP_158_296_6262/n677 ), 
	.A(\DP_OP_158_296_6262/n664 ));
   NOR2X1TS U734 (.Y(\DP_OP_158_296_6262/n630 ), 
	.B(\DP_OP_158_296_6262/n649 ), 
	.A(\DP_OP_158_296_6262/n632 ));
   NAND2X2TS U735 (.Y(\DP_OP_158_296_6262/n465 ), 
	.B(n1216), 
	.A(\DP_OP_158_296_6262/n484 ));
   NAND2X2TS U736 (.Y(\DP_OP_158_296_6262/n511 ), 
	.B(\DP_OP_158_296_6262/n549 ), 
	.A(\DP_OP_158_296_6262/n513 ));
   NAND2X1TS U737 (.Y(\DP_OP_158_296_6262/n729 ), 
	.B(\DP_OP_158_296_6262/n751 ), 
	.A(\DP_OP_158_296_6262/n731 ));
   NAND2X1TS U738 (.Y(\DP_OP_158_296_6262/n685 ), 
	.B(\DP_OP_158_296_6262/n711 ), 
	.A(\DP_OP_158_296_6262/n687 ));
   NAND2X1TS U739 (.Y(\DP_OP_158_296_6262/n628 ), 
	.B(\DP_OP_158_296_6262/n662 ), 
	.A(\DP_OP_158_296_6262/n630 ));
   NOR2X4TS U740 (.Y(\DP_OP_158_296_6262/n450 ), 
	.B(\DP_OP_158_296_6262/n452 ), 
	.A(\DP_OP_158_296_6262/n465 ));
   NOR2X4TS U741 (.Y(\DP_OP_158_296_6262/n509 ), 
	.B(\DP_OP_158_296_6262/n511 ), 
	.A(\DP_OP_158_296_6262/n576 ));
   AND2X4TS U742 (.Y(n1214), 
	.B(\DP_OP_158_296_6262/n450 ), 
	.A(\DP_OP_158_296_6262/n509 ));
   AND2X4TS U743 (.Y(n1215), 
	.B(\DP_OP_158_296_6262/n727 ), 
	.A(\DP_OP_158_296_6262/n626 ));
   NAND2X8TS U744 (.Y(\addr_calc/fft_write_calc/counter/N38 ), 
	.B(n1214), 
	.A(n1215));
   AOI21X4TS U745 (.Y(n2797), 
	.B0(FE_OFN560_n2587), 
	.A1(FE_OFN323_data_from_fft), 
	.A0(\addr_calc/fft_write_calc/counter/N38 ));
   NAND2BX1TS U746 (.Y(n1217), 
	.B(FE_OFN31_n2795), 
	.AN(n1218));
   XNOR2X1TS U747 (.Y(n1218), 
	.B(FE_OFN285_addr_calc_fft_write_calc_count_22_), 
	.A(\add_x_22_1/n34 ));
   OAI2BB1X1TS U749 (.Y(n1044), 
	.B0(n1217), 
	.A1N(FE_OFN22_n2797), 
	.A0N(FE_OFN285_addr_calc_fft_write_calc_count_22_));
   XNOR2X1TS U750 (.Y(n1221), 
	.B(FE_OFN280_addr_calc_fft_write_calc_count_20_), 
	.A(\add_x_22_1/n41 ));
   NAND2BX1TS U752 (.Y(n1220), 
	.B(FE_OFN30_n2795), 
	.AN(n1221));
   OAI2BB1X1TS U753 (.Y(n1046), 
	.B0(n1220), 
	.A1N(FE_OFN21_n2797), 
	.A0N(FE_OFN280_addr_calc_fft_write_calc_count_20_));
   CLKINVX2TS U754 (.Y(n1223), 
	.A(n1616));
   NAND2BX1TS U755 (.Y(n1226), 
	.B(\addr_calc/fir_write_calc/counter/N53 ), 
	.AN(n1758));
   OAI2BB1X1TS U756 (.Y(n1120), 
	.B0(n1226), 
	.A1N(FE_OCPUNCON1084_n2805), 
	.A0N(n1874));
   NAND2BX1TS U757 (.Y(n1225), 
	.B(\addr_calc/fir_write_calc/counter/N50 ), 
	.AN(FE_OFN47_n1758));
   OAI2BB1X1TS U758 (.Y(n1123), 
	.B0(n1225), 
	.A1N(FE_OCPUNCON1092_n2805), 
	.A0N(n1869));
   NAND2BX1TS U759 (.Y(n1224), 
	.B(\addr_calc/fir_write_calc/counter/N44 ), 
	.AN(FE_OFN47_n1758));
   OAI2BB1X1TS U760 (.Y(n1129), 
	.B0(n1224), 
	.A1N(FE_OCPUNCON1091_n2805), 
	.A0N(\addr_calc/fir_write_calc/count[1] ));
   NAND2BX1TS U761 (.Y(n1615), 
	.B(n1223), 
	.AN(FE_OFN47_n1758));
   OAI2BB1X1TS U762 (.Y(n1230), 
	.B0(n1232), 
	.A1N(n1231), 
	.A0N(FE_OFN142_add_x_19_2_n59));
   OAI2BB1X1TS U763 (.Y(n1232), 
	.B0(n1233), 
	.A1N(\add_x_19_2/n59 ), 
	.A0N(\add_x_19_2/n58 ));
   CLKINVX2TS U764 (.Y(n1233), 
	.A(n1231));
   NOR2BX1TS U765 (.Y(n1229), 
	.B(n1231), 
	.AN(FE_OFN142_add_x_19_2_n59));
   NAND2BX1TS U766 (.Y(n1227), 
	.B(n1231), 
	.AN(\add_x_19_2/n58 ));
   NOR2BX1TS U767 (.Y(n1231), 
	.B(\add_x_19_2/n55 ), 
	.AN(\add_x_19_2/n56 ));
   NOR2X8TS U768 (.Y(\DP_OP_158_296_6262/n1999 ), 
	.B(FE_OFN496_filesize_4_), 
	.A(FE_OFN495_filesize_5_));
   NOR2X6TS U769 (.Y(\DP_OP_158_296_6262/n1988 ), 
	.B(FE_OFN493_filesize_7_), 
	.A(FE_OFN494_filesize_6_));
   NAND2X8TS U770 (.Y(\DP_OP_158_296_6262/n1987 ), 
	.B(\DP_OP_158_296_6262/n1988 ), 
	.A(\DP_OP_158_296_6262/n1999 ));
   NOR2BX4TS U771 (.Y(n1234), 
	.B(FE_OFN498_filesize_3_), 
	.AN(n1641));
   NAND2X8TS U772 (.Y(\DP_OP_158_296_6262/n2011 ), 
	.B(n1797), 
	.A(n1234));
   NAND2X4TS U773 (.Y(\DP_OP_158_296_6262/n1932 ), 
	.B(\DP_OP_158_296_6262/n1933 ), 
	.A(\DP_OP_158_296_6262/n1945 ));
   NOR2X8TS U774 (.Y(\DP_OP_158_296_6262/n1931 ), 
	.B(\DP_OP_158_296_6262/n1932 ), 
	.A(\DP_OP_158_296_6262/n1958 ));
   NOR2X1TS U775 (.Y(\DP_OP_158_296_6262/n1923 ), 
	.B(FE_OFN482_filesize_16_), 
	.A(n2589));
   XNOR2X4TS U776 (.Y(n1729), 
	.B(n2369), 
	.A(\DP_OP_158_296_6262/n1923 ));
   XNOR2X1TS U777 (.Y(\DP_OP_158_296_6262/n1716 ), 
	.B(FE_OFN252_addr_calc_fir_write_calc_count_0_), 
	.A(FE_OFN518_n2372));
   XOR2X1TS U778 (.Y(n1235), 
	.B(\addr_calc/fir_write_calc/count[2] ), 
	.A(n2596));
   XOR2X1TS U779 (.Y(n1238), 
	.B(FE_OFN241_addr_calc_fir_write_calc_count_4_), 
	.A(\DP_OP_158_296_6262/n855 ));
   XOR2X1TS U780 (.Y(n1237), 
	.B(n1866), 
	.A(FE_OFN75_n2599));
   XOR2X1TS U781 (.Y(n1236), 
	.B(FE_OFN254_addr_calc_fir_write_calc_count_6_), 
	.A(n2593));
   XOR2X1TS U782 (.Y(n1239), 
	.B(\addr_calc/fir_write_calc/count[5] ), 
	.A(n2595));
   XNOR2X1TS U783 (.Y(\DP_OP_158_296_6262/n1647 ), 
	.B(n1469), 
	.A(n1872));
   XNOR2X1TS U784 (.Y(\DP_OP_158_296_6262/n1638 ), 
	.B(n1656), 
	.A(n1874));
   XNOR2X1TS U785 (.Y(\DP_OP_158_296_6262/n1607 ), 
	.B(FE_OFN524_n1659), 
	.A(n1880));
   XNOR2X1TS U786 (.Y(\DP_OP_158_296_6262/n1618 ), 
	.B(FE_OFN232_addr_calc_fir_write_calc_count_12_), 
	.A(n1756));
   XNOR2X1TS U787 (.Y(\DP_OP_158_296_6262/n1558 ), 
	.B(n1886), 
	.A(n1729));
   XNOR2X1TS U788 (.Y(\DP_OP_158_296_6262/n1543 ), 
	.B(\addr_calc/fir_write_calc/count[18] ), 
	.A(\DP_OP_158_296_6262/n841 ));
   XNOR2X1TS U789 (.Y(\DP_OP_158_296_6262/n1526 ), 
	.B(\addr_calc/fir_write_calc/count[19] ), 
	.A(n1654));
   XNOR2X2TS U790 (.Y(\DP_OP_158_296_6262/n1380 ), 
	.B(FE_OFN273_addr_calc_fir_write_calc_count_29_), 
	.A(n1463));
   XOR2X1TS U791 (.Y(\DP_OP_158_296_6262/n1460 ), 
	.B(\add_x_22_3/n22 ), 
	.A(n1718));
   XNOR2X4TS U792 (.Y(\DP_OP_158_296_6262/n1445 ), 
	.B(FE_OFN231_addr_calc_fir_write_calc_count_25_), 
	.A(n1655));
   XNOR2X1TS U793 (.Y(\DP_OP_158_296_6262/n1409 ), 
	.B(\addr_calc/fir_write_calc/count[27] ), 
	.A(n2602));
   XNOR2X4TS U794 (.Y(\DP_OP_158_296_6262/n1428 ), 
	.B(FE_OFN268_addr_calc_fir_write_calc_count_26_), 
	.A(\DP_OP_158_296_6262/n833 ));
   XOR2X1TS U795 (.Y(\DP_OP_158_296_6262/n1502 ), 
	.B(n1891), 
	.A(FE_OFN529_DP_OP_158_296_6262_n838));
   XNOR2X1TS U796 (.Y(\DP_OP_158_296_6262/n1515 ), 
	.B(FE_OFN283_addr_calc_fir_write_calc_count_20_), 
	.A(n1776));
   XNOR2X4TS U797 (.Y(\DP_OP_158_296_6262/n1474 ), 
	.B(n2563), 
	.A(n1730));
   XNOR2X4TS U798 (.Y(\DP_OP_158_296_6262/n1489 ), 
	.B(\addr_calc/fir_write_calc/count[22] ), 
	.A(n1652));
   NOR2X2TS U799 (.Y(\DP_OP_158_296_6262/n1661 ), 
	.B(\DP_OP_158_296_6262/n1670 ), 
	.A(\DP_OP_158_296_6262/n1663 ));
   NOR2X1TS U800 (.Y(\DP_OP_158_296_6262/n1645 ), 
	.B(\DP_OP_158_296_6262/n1656 ), 
	.A(\DP_OP_158_296_6262/n1647 ));
   NOR2X2TS U801 (.Y(\DP_OP_158_296_6262/n1625 ), 
	.B(\DP_OP_158_296_6262/n1627 ), 
	.A(\DP_OP_158_296_6262/n1638 ));
   NOR2X1TS U802 (.Y(\DP_OP_158_296_6262/n1581 ), 
	.B(\DP_OP_158_296_6262/n1583 ), 
	.A(\DP_OP_158_296_6262/n1596 ));
   NOR2X1TS U803 (.Y(\DP_OP_158_296_6262/n1605 ), 
	.B(\DP_OP_158_296_6262/n1607 ), 
	.A(\DP_OP_158_296_6262/n1618 ));
   NOR2X1TS U804 (.Y(\DP_OP_158_296_6262/n1556 ), 
	.B(\DP_OP_158_296_6262/n1571 ), 
	.A(\DP_OP_158_296_6262/n1558 ));
   NOR2X2TS U805 (.Y(\DP_OP_158_296_6262/n1524 ), 
	.B(\DP_OP_158_296_6262/n1543 ), 
	.A(\DP_OP_158_296_6262/n1526 ));
   XOR2X4TS U806 (.Y(n1240), 
	.B(FE_OFN238_addr_calc_fir_write_calc_count_30_), 
	.A(\DP_OP_158_296_6262/n829 ));
   NOR2X4TS U807 (.Y(\DP_OP_158_296_6262/n1378 ), 
	.B(\DP_OP_158_296_6262/n1395 ), 
	.A(\DP_OP_158_296_6262/n1380 ));
   NOR2X1TS U808 (.Y(\DP_OP_158_296_6262/n1443 ), 
	.B(\DP_OP_158_296_6262/n1460 ), 
	.A(\DP_OP_158_296_6262/n1445 ));
   NOR2X2TS U809 (.Y(\DP_OP_158_296_6262/n1407 ), 
	.B(\DP_OP_158_296_6262/n1409 ), 
	.A(\DP_OP_158_296_6262/n1428 ));
   NOR2X1TS U810 (.Y(\DP_OP_158_296_6262/n1500 ), 
	.B(\DP_OP_158_296_6262/n1502 ), 
	.A(\DP_OP_158_296_6262/n1515 ));
   NOR2X2TS U811 (.Y(\DP_OP_158_296_6262/n1472 ), 
	.B(\DP_OP_158_296_6262/n1489 ), 
	.A(\DP_OP_158_296_6262/n1474 ));
   NAND2X2TS U812 (.Y(\DP_OP_158_296_6262/n1659 ), 
	.B(\DP_OP_158_296_6262/n1688 ), 
	.A(\DP_OP_158_296_6262/n1661 ));
   NAND2X1TS U813 (.Y(\DP_OP_158_296_6262/n1623 ), 
	.B(\DP_OP_158_296_6262/n1645 ), 
	.A(\DP_OP_158_296_6262/n1625 ));
   NAND2X2TS U814 (.Y(\DP_OP_158_296_6262/n1579 ), 
	.B(\DP_OP_158_296_6262/n1581 ), 
	.A(\DP_OP_158_296_6262/n1605 ));
   NAND2X2TS U815 (.Y(\DP_OP_158_296_6262/n1522 ), 
	.B(\DP_OP_158_296_6262/n1556 ), 
	.A(\DP_OP_158_296_6262/n1524 ));
   NAND2X4TS U816 (.Y(\DP_OP_158_296_6262/n1359 ), 
	.B(n1240), 
	.A(\DP_OP_158_296_6262/n1378 ));
   NAND2X1TS U817 (.Y(\DP_OP_158_296_6262/n1405 ), 
	.B(\DP_OP_158_296_6262/n1443 ), 
	.A(\DP_OP_158_296_6262/n1407 ));
   NAND2X2TS U818 (.Y(\DP_OP_158_296_6262/n1470 ), 
	.B(\DP_OP_158_296_6262/n1500 ), 
	.A(\DP_OP_158_296_6262/n1472 ));
   NOR2X2TS U819 (.Y(\DP_OP_158_296_6262/n1621 ), 
	.B(FE_OFN538_DP_OP_158_296_6262_n1659), 
	.A(\DP_OP_158_296_6262/n1623 ));
   NOR2X4TS U820 (.Y(\DP_OP_158_296_6262/n1520 ), 
	.B(\DP_OP_158_296_6262/n1579 ), 
	.A(\DP_OP_158_296_6262/n1522 ));
   NOR2X4TS U821 (.Y(\DP_OP_158_296_6262/n1344 ), 
	.B(\DP_OP_158_296_6262/n1346 ), 
	.A(\DP_OP_158_296_6262/n1359 ));
   NOR2X4TS U822 (.Y(\DP_OP_158_296_6262/n1403 ), 
	.B(\DP_OP_158_296_6262/n1405 ), 
	.A(\DP_OP_158_296_6262/n1470 ));
   NAND2X4TS U823 (.Y(\DP_OP_158_296_6262/n1518 ), 
	.B(\DP_OP_158_296_6262/n1621 ), 
	.A(\DP_OP_158_296_6262/n1520 ));
   NAND2X6TS U824 (.Y(\DP_OP_158_296_6262/n1342 ), 
	.B(\DP_OP_158_296_6262/n1344 ), 
	.A(\DP_OP_158_296_6262/n1403 ));
   OR2X8TS U825 (.Y(\addr_calc/fir_write_calc/counter/N38 ), 
	.B(\DP_OP_158_296_6262/n1518 ), 
	.A(\DP_OP_158_296_6262/n1342 ));
   OR3X1TS U826 (.Y(n1241), 
	.C(n2061), 
	.B(n2804), 
	.A(FE_OFN318_data_cntl_N95));
   CLKINVX1TS U827 (.Y(\add_x_22_3/n121 ), 
	.A(\addr_calc/fir_write_calc/count[1] ));
   XNOR2X1TS U828 (.Y(\addr_calc/fir_write_calc/counter/N44 ), 
	.B(\addr_calc/fir_write_calc/count[0] ), 
	.A(\add_x_22_3/n121 ));
   XNOR2X1TS U829 (.Y(n1243), 
	.B(\addr_calc/fft_write_calc/count[6] ), 
	.A(\add_x_22_1/n102 ));
   NAND2BX1TS U831 (.Y(n1242), 
	.B(FE_OFN35_n2795), 
	.AN(n1243));
   OAI2BB1X1TS U832 (.Y(n1060), 
	.B0(n1242), 
	.A1N(FE_OFN26_n2797), 
	.A0N(\addr_calc/fft_write_calc/count[6] ));
   NAND2X4TS U833 (.Y(\DP_OP_159_297_3515/n1039 ), 
	.B(\DP_OP_159_297_3515/n1040 ), 
	.A(\DP_OP_159_297_3515/n1064 ));
   NOR2X1TS U834 (.Y(\DP_OP_159_297_3515/n985 ), 
	.B(\DP_OP_159_297_3515/n986 ), 
	.A(\DP_OP_159_297_3515/n998 ));
   AND2X4TS U835 (.Y(n1245), 
	.B(\DP_OP_159_297_3515/n1011 ), 
	.A(\DP_OP_159_297_3515/n985 ));
   NAND2BX4TS U836 (.Y(n1782), 
	.B(n1245), 
	.AN(FE_OFN519_DP_OP_159_297_3515_n1039));
   CLKINVX1TS U837 (.Y(\DP_OP_159_297_3515/n970 ), 
	.A(\DP_OP_159_297_3515/n971 ));
   NAND2X1TS U838 (.Y(\DP_OP_159_297_3515/n969 ), 
	.B(\DP_OP_159_297_3515/n970 ), 
	.A(FE_OFN553_n1789));
   XNOR2X4TS U839 (.Y(n1662), 
	.B(\DP_OP_159_297_3515/n964 ), 
	.A(\DP_OP_159_297_3515/n969 ));
   XNOR2X1TS U840 (.Y(\DP_OP_159_297_3515/n353 ), 
	.B(\DP_OP_159_297_3515/n815 ), 
	.A(\addr_calc/iir_read_calc/count[0] ));
   XOR2X1TS U841 (.Y(n1246), 
	.B(\addr_calc/iir_read_calc/count[2] ), 
	.A(n2612));
   XOR2X1TS U842 (.Y(n1248), 
	.B(FE_OFN244_addr_calc_iir_read_calc_count_4_), 
	.A(n2624));
   NOR2X1TS U843 (.Y(\DP_OP_159_297_3515/n339 ), 
	.B(\DP_OP_159_297_3515/n341 ), 
	.A(\DP_OP_159_297_3515/n343 ));
   XOR2X1TS U844 (.Y(n1249), 
	.B(n2553), 
	.A(n2623));
   XOR2X1TS U845 (.Y(n1247), 
	.B(n2018), 
	.A(n2610));
   NAND2X1TS U846 (.Y(\DP_OP_159_297_3515/n333 ), 
	.B(n1248), 
	.A(\DP_OP_159_297_3515/n339 ));
   XNOR2X1TS U847 (.Y(\DP_OP_159_297_3515/n305 ), 
	.B(n2583), 
	.A(n2622));
   XNOR2X1TS U848 (.Y(\DP_OP_159_297_3515/n298 ), 
	.B(\addr_calc/iir_read_calc/count[9] ), 
	.A(n2608));
   XNOR2X1TS U849 (.Y(\DP_OP_159_297_3515/n280 ), 
	.B(FE_OFN236_addr_calc_iir_read_calc_count_11_), 
	.A(n2620));
   XOR2X1TS U850 (.Y(\DP_OP_159_297_3515/n260 ), 
	.B(\add_x_22_4/n71 ), 
	.A(n2618));
   XNOR2X1TS U851 (.Y(\DP_OP_159_297_3515/n249 ), 
	.B(n1784), 
	.A(n2617));
   XNOR2X1TS U852 (.Y(\DP_OP_159_297_3515/n225 ), 
	.B(n1916), 
	.A(n2615));
   XNOR2X1TS U853 (.Y(\DP_OP_159_297_3515/n238 ), 
	.B(n2566), 
	.A(n2616));
   XNOR2X2TS U854 (.Y(\DP_OP_159_297_3515/n200 ), 
	.B(n2024), 
	.A(\DP_OP_159_297_3515/n1128 ));
   XNOR2X1TS U855 (.Y(\DP_OP_159_297_3515/n213 ), 
	.B(\addr_calc/iir_read_calc/count[17] ), 
	.A(n2607));
   XNOR2X4TS U856 (.Y(\DP_OP_159_297_3515/n185 ), 
	.B(n2556), 
	.A(n1662));
   XOR2X4TS U857 (.Y(\DP_OP_159_297_3515/n168 ), 
	.B(n2027), 
	.A(n1697));
   NOR2X2TS U858 (.Y(\DP_OP_159_297_3515/n315 ), 
	.B(\DP_OP_159_297_3515/n333 ), 
	.A(\DP_OP_159_297_3515/n317 ));
   NOR2X1TS U859 (.Y(\DP_OP_159_297_3515/n303 ), 
	.B(\DP_OP_159_297_3515/n312 ), 
	.A(\DP_OP_159_297_3515/n305 ));
   NOR2X1TS U860 (.Y(\DP_OP_159_297_3515/n287 ), 
	.B(\DP_OP_159_297_3515/n298 ), 
	.A(\DP_OP_159_297_3515/n289 ));
   NOR2X1TS U861 (.Y(\DP_OP_159_297_3515/n267 ), 
	.B(\DP_OP_159_297_3515/n269 ), 
	.A(\DP_OP_159_297_3515/n280 ));
   NOR2X1TS U862 (.Y(\DP_OP_159_297_3515/n247 ), 
	.B(\DP_OP_159_297_3515/n260 ), 
	.A(\DP_OP_159_297_3515/n249 ));
   NOR2X1TS U863 (.Y(\DP_OP_159_297_3515/n223 ), 
	.B(\DP_OP_159_297_3515/n225 ), 
	.A(\DP_OP_159_297_3515/n238 ));
   NOR2X2TS U864 (.Y(\DP_OP_159_297_3515/n198 ), 
	.B(\DP_OP_159_297_3515/n200 ), 
	.A(\DP_OP_159_297_3515/n213 ));
   NOR2X2TS U865 (.Y(\DP_OP_159_297_3515/n166 ), 
	.B(\DP_OP_159_297_3515/n185 ), 
	.A(\DP_OP_159_297_3515/n168 ));
   NAND2X2TS U866 (.Y(\DP_OP_159_297_3515/n301 ), 
	.B(\DP_OP_159_297_3515/n315 ), 
	.A(\DP_OP_159_297_3515/n303 ));
   NAND2X1TS U867 (.Y(\DP_OP_159_297_3515/n265 ), 
	.B(\DP_OP_159_297_3515/n287 ), 
	.A(\DP_OP_159_297_3515/n267 ));
   NAND2X1TS U868 (.Y(\DP_OP_159_297_3515/n221 ), 
	.B(\DP_OP_159_297_3515/n247 ), 
	.A(\DP_OP_159_297_3515/n223 ));
   NAND2X4TS U869 (.Y(\DP_OP_159_297_3515/n164 ), 
	.B(\DP_OP_159_297_3515/n198 ), 
	.A(\DP_OP_159_297_3515/n166 ));
   NOR2X2TS U870 (.Y(\DP_OP_159_297_3515/n263 ), 
	.B(FE_OFN537_DP_OP_159_297_3515_n301), 
	.A(\DP_OP_159_297_3515/n265 ));
   NOR2X4TS U871 (.Y(\DP_OP_159_297_3515/n162 ), 
	.B(\DP_OP_159_297_3515/n221 ), 
	.A(\DP_OP_159_297_3515/n164 ));
   NAND2X4TS U872 (.Y(\DP_OP_159_297_3515/n160 ), 
	.B(\DP_OP_159_297_3515/n263 ), 
	.A(\DP_OP_159_297_3515/n162 ));
   OR2X2TS U873 (.Y(\addr_calc/iir_read_calc/counter/N38 ), 
	.B(\DP_OP_159_297_3515/n160 ), 
	.A(\DP_OP_159_297_3515/n1 ));
   OAI21XLTS U874 (.Y(n1250), 
	.B0(iir_enable), 
	.A1(n2785), 
	.A0(n2786));
   XNOR2X1TS U875 (.Y(n1253), 
	.B(\add_x_22_4/n71 ), 
	.A(n1254));
   NAND2BX1TS U876 (.Y(n1254), 
	.B(\add_x_22_4/n75 ), 
	.AN(n1255));
   CLKINVX2TS U877 (.Y(n1255), 
	.A(n1785));
   CLKINVX2TS U878 (.Y(n1251), 
	.A(\add_x_22_4/n71 ));
   NAND2BX1TS U879 (.Y(n1252), 
	.B(FE_OCPUNCON1878_n2787), 
	.AN(n1253));
   OAI2BB1X1TS U880 (.Y(n958), 
	.B0(n1252), 
	.A1N(FE_OFN85_n2654), 
	.A0N(n1251));
   NOR2X1TS U881 (.Y(\DP_OP_158_296_6262/n1174 ), 
	.B(\DP_OP_158_296_6262/n1212 ), 
	.A(\DP_OP_158_296_6262/n1176 ));
   OAI2BB1X1TS U897 (.Y(n1126), 
	.B0(n1615), 
	.A1N(FE_OCPUNCON1092_n2805), 
	.A0N(\addr_calc/fir_write_calc/count[4] ));
   XOR2X4TS U898 (.Y(n1623), 
	.B(FE_OFN286_addr_calc_iir_read_calc_count_30_), 
	.A(n2625));
   XNOR2X1TS U899 (.Y(\DP_OP_159_297_3515/n430 ), 
	.B(\addr_calc/iir_write_calc/count[31] ), 
	.A(n2614));
   INVX2TS U900 (.Y(n1733), 
	.A(\DP_OP_159_297_3515/n1024 ));
   XNOR2X1TS U901 (.Y(n1563), 
	.B(n1850), 
	.A(n2613));
   CLKXOR2X4TS U902 (.Y(n2598), 
	.B(n2364), 
	.A(n1693));
   NOR2X2TS U903 (.Y(\add_x_19_5/n118 ), 
	.B(\add_x_19_5/n120 ), 
	.A(\add_x_19_5/n123 ));
   NOR2X4TS U904 (.Y(\add_x_19_0/n55 ), 
	.B(FE_OFN356_offset_27_), 
	.A(n1944));
   NOR2X4TS U905 (.Y(\add_x_19_5/n55 ), 
	.B(FE_OFN355_offset_27_), 
	.A(n1688));
   NOR2X1TS U907 (.Y(\add_x_19_2/n86 ), 
	.B(FE_OCPUNCON1070_FE_OFN377_offset_21_), 
	.A(n1879));
   NOR2X1TS U908 (.Y(n1555), 
	.B(n1557), 
	.A(n1556));
   NOR2X1TS U909 (.Y(n1557), 
	.B(FE_OFN338_offset_31_), 
	.A(FE_OFN274_addr_calc_fft_write_calc_count_31_));
   AND2X2TS U910 (.Y(n1556), 
	.B(FE_OFN338_offset_31_), 
	.A(FE_OFN274_addr_calc_fft_write_calc_count_31_));
   NOR2BX1TS U911 (.Y(n1552), 
	.B(n1555), 
	.AN(\add_x_19_1/n37 ));
   INVX2TS U912 (.Y(n1554), 
	.A(n1555));
   INVX2TS U913 (.Y(n1546), 
	.A(\add_x_19_1/n42 ));
   NOR2BX1TS U914 (.Y(n1575), 
	.B(\add_x_22_5/n67 ), 
	.AN(\add_x_22_5/n68 ));
   NOR2BX1TS U915 (.Y(n1578), 
	.B(\add_x_22_4/n15 ), 
	.AN(\add_x_22_4/n16 ));
   NOR2BX1TS U916 (.Y(n1622), 
	.B(\add_x_22_0/n85 ), 
	.AN(n1972));
   INVX2TS U918 (.Y(n1572), 
	.A(\add_x_22_4/n15 ));
   INVX2TS U920 (.Y(n1541), 
	.A(\add_x_19_0/n42 ));
   NOR2X2TS U921 (.Y(\add_x_19_3/n55 ), 
	.B(FE_OFN356_offset_27_), 
	.A(n1835));
   NOR2BX1TS U923 (.Y(n1605), 
	.B(n1607), 
	.AN(FE_OFN144_add_x_19_5_n59));
   NOR2BX1TS U924 (.Y(n1607), 
	.B(\add_x_19_5/n55 ), 
	.AN(\add_x_19_5/n56 ));
   NOR2BX1TS U925 (.Y(n1635), 
	.B(\add_x_22_0/n58 ), 
	.AN(n2554));
   NAND2BX1TS U926 (.Y(n1629), 
	.B(\add_x_22_0/n41 ), 
	.AN(\add_x_22_0/n40 ));
   INVX2TS U928 (.Y(\add_x_22_4/n15 ), 
	.A(\addr_calc/iir_read_calc/count[26] ));
   XNOR2X1TS U929 (.Y(n2599), 
	.B(FE_OFN498_filesize_3_), 
	.A(\DP_OP_158_296_6262/n2015 ));
   NOR2X2TS U930 (.Y(\add_x_19_2/n118 ), 
	.B(\add_x_19_2/n120 ), 
	.A(\add_x_19_2/n123 ));
   XNOR2X1TS U931 (.Y(\DP_OP_158_296_6262/n161 ), 
	.B(\addr_calc/fir_read_calc/count[21] ), 
	.A(FE_OFN529_DP_OP_158_296_6262_n838));
   NOR2BX1TS U932 (.Y(n1625), 
	.B(n2796), 
	.AN(n1626));
   NOR2X1TS U933 (.Y(n1626), 
	.B(FE_OFN322_data_cntl_N9), 
	.A(FE_OFN560_n2587));
   OAI21X4TS U934 (.Y(n1595), 
	.B0(\add_x_19_3/n121 ), 
	.A1(\add_x_19_3/n124 ), 
	.A0(\add_x_19_3/n120 ));
   NOR2X4TS U935 (.Y(n1558), 
	.B(\add_x_19_0/n165 ), 
	.A(\add_x_19_0/n162 ));
   CLKINVX2TS U936 (.Y(\DP_OP_158_296_6262/n1897 ), 
	.A(FE_OFN477_filesize_20_));
   NOR2X1TS U937 (.Y(\add_x_19_4/n63 ), 
	.B(FE_OFN364_offset_25_), 
	.A(n1926));
   NOR2X4TS U938 (.Y(\add_x_19_0/n78 ), 
	.B(FE_OFN371_offset_23_), 
	.A(n1950));
   OAI21X2TS U939 (.Y(\add_x_19_0/n85 ), 
	.B0(\add_x_19_0/n87 ), 
	.A1(\add_x_19_0/n86 ), 
	.A0(\add_x_19_0/n90 ));
   NOR2X2TS U940 (.Y(\DP_OP_158_296_6262/n304 ), 
	.B(\DP_OP_158_296_6262/n315 ), 
	.A(\DP_OP_158_296_6262/n306 ));
   NOR2X2TS U941 (.Y(\add_x_19_0/n120 ), 
	.B(FE_OFN400_offset_15_), 
	.A(n1689));
   NOR2X4TS U942 (.Y(\add_x_19_5/n78 ), 
	.B(FE_OFN372_offset_23_), 
	.A(n1965));
   NOR4XLTS U943 (.Y(n918), 
	.D(n1974), 
	.C(\addr_calc/iir_write_calc/count[29] ), 
	.B(n2036), 
	.A(FE_OFN239_addr_calc_iir_write_calc_count_30_));
   NOR2X1TS U944 (.Y(\add_x_19_4/n61 ), 
	.B(\add_x_19_4/n63 ), 
	.A(\add_x_19_4/n66 ));
   NOR2X1TS U945 (.Y(\add_x_19_1/n55 ), 
	.B(FE_OFN353_offset_27_), 
	.A(n1913));
   NOR2X1TS U947 (.Y(\add_x_19_1/n139 ), 
	.B(FE_OCPN1905_FE_OCPUNCON1873_offset_11_), 
	.A(n1667));
   NOR2X2TS U948 (.Y(\add_x_19_5/n114 ), 
	.B(\add_x_19_5/n116 ), 
	.A(\add_x_19_5/n135 ));
   NOR2X1TS U949 (.Y(\add_x_19_2/n48 ), 
	.B(n1871), 
	.A(FE_OFN350_offset_28_));
   OAI21X4TS U950 (.Y(n1588), 
	.B0(\add_x_19_0/n182 ), 
	.A1(\add_x_19_0/n185 ), 
	.A0(\add_x_19_0/n181 ));
   OAI21X2TS U952 (.Y(\add_x_19_1/n187 ), 
	.B0(\add_x_19_1/n189 ), 
	.A1(\add_x_19_1/n191 ), 
	.A0(\add_x_19_1/n188 ));
   INVX2TS U953 (.Y(n2066), 
	.A(n2065));
   NOR2X1TS U956 (.Y(\add_x_19_1/n123 ), 
	.B(FE_OFN403_offset_14_), 
	.A(FE_OFN259_addr_calc_fft_write_calc_count_14_));
   NOR2X4TS U957 (.Y(\add_x_19_5/n97 ), 
	.B(FE_OFN384_offset_19_), 
	.A(n1958));
   INVXLTS U958 (.Y(\add_x_22_4/n67 ), 
	.A(\addr_calc/iir_read_calc/count[14] ));
   INVX2TS U959 (.Y(\add_x_22_4/n74 ), 
	.A(\addr_calc/iir_read_calc/count[12] ));
   OAI2BB1X1TS U964 (.Y(n1534), 
	.B0(\add_x_19_5/n37 ), 
	.A1N(n1589), 
	.A0N(n1533));
   NOR2BX1TS U965 (.Y(n1532), 
	.B(\add_x_19_5/n36 ), 
	.AN(n2629));
   NOR2BX1TS U967 (.Y(n1640), 
	.B(\add_x_19_4/n36 ), 
	.AN(\add_x_19_4/n37 ));
   INVX2TS U968 (.Y(n1583), 
	.A(\add_x_19_4/n40 ));
   OA21XLTS U969 (.Y(n1585), 
	.B0(\add_x_19_4/n37 ), 
	.A1(n1583), 
	.A0(\add_x_19_4/n36 ));
   NOR2BX1TS U970 (.Y(n1584), 
	.B(\add_x_19_4/n36 ), 
	.AN(n2634));
   INVX2TS U971 (.Y(n1589), 
	.A(\add_x_19_5/n42 ));
   NOR2X2TS U975 (.Y(n2793), 
	.B(n1298), 
	.A(n1297));
   INVX2TS U977 (.Y(n2005), 
	.A(\addr_calc/fir_write_calc/count[18] ));
   INVX2TS U979 (.Y(n1878), 
	.A(\addr_calc/fir_read_calc/count[21] ));
   NOR2X4TS U982 (.Y(\add_x_19_4/n170 ), 
	.B(\addr_calc/iir_read_calc/count[5] ), 
	.A(FE_OCP_RBN1492_offset_5_));
   NAND2X1TS U983 (.Y(\add_x_19_4/n124 ), 
	.B(\addr_calc/iir_read_calc/count[14] ), 
	.A(FE_OFN405_offset_14_));
   NAND2X4TS U984 (.Y(\add_x_19_3/n132 ), 
	.B(FE_OFN413_offset_12_), 
	.A(FE_OFN232_addr_calc_fir_write_calc_count_12_));
   NOR2X1TS U985 (.Y(\add_x_19_2/n123 ), 
	.B(FE_OFN402_offset_14_), 
	.A(n1690));
   NAND2X1TS U986 (.Y(\add_x_19_1/n67 ), 
	.B(FE_OFN365_offset_24_), 
	.A(FE_OFN277_addr_calc_fft_write_calc_count_24_));
   NOR2X1TS U987 (.Y(\add_x_19_0/n123 ), 
	.B(FE_OFN404_offset_14_), 
	.A(n2043));
   NAND2X8TS U988 (.Y(\add_x_19_5/n111 ), 
	.B(\addr_calc/iir_write_calc/count[16] ), 
	.A(FE_OFN397_offset_16_));
   NAND2X2TS U990 (.Y(\add_x_19_3/n155 ), 
	.B(FE_OFN255_addr_calc_fir_write_calc_count_8_), 
	.A(FE_OFN428_offset_8_));
   NOR2X2TS U991 (.Y(\add_x_19_1/n165 ), 
	.B(FE_OCPUNCON1684_offset_6_), 
	.A(FE_OFN271_addr_calc_fft_write_calc_count_6_));
   NOR2X8TS U992 (.Y(\add_x_19_0/n162 ), 
	.B(n1666), 
	.A(FE_OCPUNCON1278_offset_7_));
   NOR2X4TS U993 (.Y(\add_x_19_4/n181 ), 
	.B(FE_OCPUNCON1075_FE_OFN447_offset_3_), 
	.A(n1902));
   INVX2TS U994 (.Y(n2060), 
	.A(FE_OFN565_n2066));
   INVX8TS U995 (.Y(\DP_OP_158_296_6262/n829 ), 
	.A(\DP_OP_158_296_6262/n2060 ));
   INVX2TS U996 (.Y(n1861), 
	.A(n2063));
   INVX2TS U997 (.Y(n2588), 
	.A(n2074));
   CLKXOR2X2TS U999 (.Y(n2596), 
	.B(n1680), 
	.A(\DP_OP_158_296_6262/n2020 ));
   CLKINVX12TS U1000 (.Y(n1718), 
	.A(\DP_OP_158_296_6262/n2054 ));
   INVX6TS U1001 (.Y(\DP_OP_158_296_6262/n833 ), 
	.A(\DP_OP_158_296_6262/n2056 ));
   INVX2TS U1002 (.Y(n1667), 
	.A(n1930));
   INVX2TS U1004 (.Y(\DP_OP_159_297_3515/n880 ), 
	.A(FE_OFN496_filesize_4_));
   NAND2BX1TS U1005 (.Y(n1569), 
	.B(\add_x_19_2/n87 ), 
	.AN(\add_x_19_2/n86 ));
   NAND2BX1TS U1006 (.Y(n1550), 
	.B(n1555), 
	.AN(\add_x_19_1/n36 ));
   AOI2BB2X1TS U1007 (.Y(n1553), 
	.B1(\add_x_19_1/n36 ), 
	.B0(n1552), 
	.A1N(n1554), 
	.A0N(\add_x_19_1/n37 ));
   XNOR2X2TS U1008 (.Y(\addr_calc/fft_write_addr[21] ), 
	.B(\add_x_19_1/n11 ), 
	.A(\add_x_19_1/n88 ));
   NAND2BX1TS U1009 (.Y(n1542), 
	.B(FE_OFN4_n1755), 
	.AN(n1543));
   NAND2BX1TS U1010 (.Y(n1565), 
	.B(FE_OCPUNCON1881_n2813), 
	.AN(n1566));
   XNOR2X1TS U1011 (.Y(n1566), 
	.B(\add_x_22_5/n57 ), 
	.A(\add_x_22_5/n58 ));
   XNOR2X1TS U1012 (.Y(n1574), 
	.B(\addr_calc/iir_write_calc/count[15] ), 
	.A(n1575));
   XNOR2X1TS U1013 (.Y(n1647), 
	.B(FE_OFN233_addr_calc_fir_write_calc_count_12_), 
	.A(\add_x_22_3/n75 ));
   XNOR2X1TS U1014 (.Y(n1577), 
	.B(\addr_calc/iir_read_calc/count[27] ), 
	.A(n1578));
   NAND2BX2TS U1015 (.Y(n1597), 
	.B(\add_x_19_2/n79 ), 
	.AN(\add_x_19_2/n78 ));
   XNOR2X1TS U1016 (.Y(n1616), 
	.B(\add_x_22_3/n109 ), 
	.A(\add_x_22_3/n110 ));
   OAI2BB2XLTS U1017 (.Y(n991), 
	.B1(\add_x_22_5/n80 ), 
	.B0(n1740), 
	.A1N(\addr_calc/iir_write_calc/counter/N54 ), 
	.A0N(FE_OCPUNCON1879_n2813));
   NAND2X1TS U1018 (.Y(n1620), 
	.B(n1621), 
	.A(n1754));
   XNOR2X1TS U1019 (.Y(n1621), 
	.B(\add_x_22_0/n80 ), 
	.A(n1622));
   XNOR2X1TS U1020 (.Y(n1609), 
	.B(FE_OFN224_addr_calc_fft_read_calc_count_6_), 
	.A(\add_x_22_0/n102 ));
   XNOR2X1TS U1021 (.Y(n1644), 
	.B(\add_x_22_0/n109 ), 
	.A(\add_x_22_0/n110 ));
   XNOR2X1TS U1022 (.Y(n1639), 
	.B(\add_x_22_0/n57 ), 
	.A(\add_x_22_0/n58 ));
   XNOR2X1TS U1023 (.Y(n1637), 
	.B(n2569), 
	.A(\add_x_22_0/n50 ));
   XNOR2X1TS U1024 (.Y(n1631), 
	.B(n2575), 
	.A(\add_x_22_0/n16 ));
   XNOR2X1TS U1025 (.Y(n1571), 
	.B(n1572), 
	.A(\add_x_22_4/n16 ));
   OAI2BB1XLTS U1026 (.Y(n1072), 
	.B0(n1612), 
	.A1N(FE_OFN69_n2809), 
	.A0N(\addr_calc/fir_read_calc/count[26] ));
   XNOR2X1TS U1027 (.Y(n1613), 
	.B(\addr_calc/fir_read_calc/count[26] ), 
	.A(\add_x_22_2/n16 ));
   NAND2BX1TS U1029 (.Y(n1537), 
	.B(\add_x_19_5/n121 ), 
	.AN(\add_x_19_5/n120 ));
   NOR2BX1TS U1030 (.Y(n1544), 
	.B(\add_x_19_0/n36 ), 
	.AN(\add_x_19_0/n37 ));
   NOR2BX1TS U1031 (.Y(n1538), 
	.B(\add_x_19_3/n36 ), 
	.AN(\add_x_19_3/n37 ));
   NAND2BX1TS U1032 (.Y(n1603), 
	.B(n1607), 
	.AN(\add_x_19_5/n58 ));
   XNOR2X1TS U1033 (.Y(n1619), 
	.B(FE_OFN282_addr_calc_fir_write_calc_count_20_), 
	.A(\add_x_22_3/n41 ));
   NAND2X1TS U1034 (.Y(n1627), 
	.B(n1628), 
	.A(FE_OFN2_n1754));
   XNOR2X1TS U1035 (.Y(n1628), 
	.B(\addr_calc/fft_read_calc/count[21] ), 
	.A(n1629));
   XNOR2X1TS U1036 (.Y(\DP_OP_158_296_6262/n1149 ), 
	.B(n2043), 
	.A(n1657));
   XNOR2X1TS U1037 (.Y(\DP_OP_158_296_6262/n1055 ), 
	.B(FE_OFN288_addr_calc_fft_read_calc_count_21_), 
	.A(FE_OFN529_DP_OP_158_296_6262_n838));
   XNOR2X1TS U1038 (.Y(\DP_OP_158_296_6262/n1124 ), 
	.B(\addr_calc/fft_read_calc/count[16] ), 
	.A(n2594));
   XNOR2X4TS U1039 (.Y(n2614), 
	.B(n2324), 
	.A(\DP_OP_159_297_3515/n885 ));
   XNOR2X2TS U1040 (.Y(n2622), 
	.B(\DP_OP_159_297_3515/n876 ), 
	.A(\DP_OP_159_297_3515/n1044 ));
   XNOR2X2TS U1041 (.Y(n1624), 
	.B(n1839), 
	.A(n2613));
   NOR2X1TS U1043 (.Y(\DP_OP_159_297_3515/n990 ), 
	.B(\DP_OP_159_297_3515/n991 ), 
	.A(\DP_OP_159_297_3515/n1012 ));
   NOR2X1TS U1044 (.Y(\DP_OP_158_296_6262/n2015 ), 
	.B(n1680), 
	.A(\DP_OP_158_296_6262/n2020 ));
   NAND2X2TS U1045 (.Y(\DP_OP_158_296_6262/n1841 ), 
	.B(\DP_OP_158_296_6262/n1842 ), 
	.A(FE_OFN113_DP_OP_158_296_6262_n1791));
   NOR2X1TS U1046 (.Y(\DP_OP_158_296_6262/n1938 ), 
	.B(FE_OFN486_filesize_14_), 
	.A(\DP_OP_158_296_6262/n1946 ));
   CLKINVX2TS U1047 (.Y(n2343), 
	.A(FE_OFN468_filesize_26_));
   INVX2TS U1048 (.Y(n1464), 
	.A(FE_OFN465_filesize_29_));
   INVX2TS U1050 (.Y(\DP_OP_159_297_3515/n792 ), 
	.A(\DP_OP_159_297_3515/n1133 ));
   NOR2X2TS U1055 (.Y(\add_x_22_3/n59 ), 
	.B(n1273), 
	.A(\add_x_22_3/n94 ));
   NAND4BX1TS U1056 (.Y(n1274), 
	.D(\add_x_22_0/n77 ), 
	.C(n1689), 
	.B(n2043), 
	.AN(\add_x_22_0/n69 ));
   NOR2X2TS U1057 (.Y(\add_x_22_0/n59 ), 
	.B(n1274), 
	.A(\add_x_22_0/n94 ));
   NAND3X1TS U1058 (.Y(n1275), 
	.C(\add_x_22_4/n77 ), 
	.B(\addr_calc/iir_read_calc/count[14] ), 
	.A(\addr_calc/iir_read_calc/count[15] ));
   NOR3X1TS U1059 (.Y(\add_x_22_4/n59 ), 
	.C(n1275), 
	.B(\add_x_22_4/n69 ), 
	.A(\add_x_22_4/n94 ));
   NAND3X1TS U1060 (.Y(n1276), 
	.C(\add_x_22_2/n77 ), 
	.B(n1690), 
	.A(n1890));
   NOR3X1TS U1061 (.Y(\add_x_22_2/n59 ), 
	.C(n1276), 
	.B(\add_x_22_2/n69 ), 
	.A(\add_x_22_2/n94 ));
   NAND2BX1TS U1062 (.Y(n1277), 
	.B(\add_x_19_2/n37 ), 
	.AN(\add_x_19_2/n36 ));
   NAND2BX1TS U1064 (.Y(n1278), 
	.B(\add_x_19_0/n67 ), 
	.AN(\add_x_19_0/n66 ));
   XOR2X4TS U1065 (.Y(\addr_calc/fft_read_addr[24] ), 
	.B(n1278), 
	.A(\add_x_19_0/n68 ));
   NAND2BX1TS U1066 (.Y(n1279), 
	.B(\add_x_19_4/n90 ), 
	.AN(\add_x_19_4/n89 ));
   NAND2BX1TS U1068 (.Y(n1280), 
	.B(\add_x_19_2/n166 ), 
	.AN(\add_x_19_2/n165 ));
   XOR2X1TS U1069 (.Y(\addr_calc/fir_read_addr[6] ), 
	.B(n1280), 
	.A(\add_x_19_2/n167 ));
   NAND2BX1TS U1070 (.Y(n1281), 
	.B(\add_x_19_1/n166 ), 
	.AN(\add_x_19_1/n165 ));
   XOR2X1TS U1071 (.Y(\addr_calc/fft_write_addr[6] ), 
	.B(n1281), 
	.A(\add_x_19_1/n167 ));
   OAI21X1TS U1072 (.Y(n1282), 
	.B0(\add_x_19_3/n155 ), 
	.A1(\add_x_19_3/n156 ), 
	.A0(\add_x_19_3/n154 ));
   CLKINVX1TS U1073 (.Y(n1283), 
	.A(\add_x_19_3/n152 ));
   OAI21X1TS U1076 (.Y(n1285), 
	.B0(\add_x_19_4/n185 ), 
	.A1(\add_x_19_4/n186 ), 
	.A0(\add_x_19_4/n184 ));
   CLKINVX1TS U1077 (.Y(n1286), 
	.A(\add_x_19_4/n182 ));
   OAI21X1TS U1078 (.Y(n1287), 
	.B0(n1285), 
	.A1(n1286), 
	.A0(\add_x_19_4/n181 ));
   OAI31X1TS U1079 (.Y(\addr_calc/iir_read_addr[3] ), 
	.B0(n1287), 
	.A2(n1286), 
	.A1(n1285), 
	.A0(\add_x_19_4/n181 ));
   OA21XLTS U1080 (.Y(\addr_calc/iir_write_addr[0] ), 
	.B0(\add_x_19_5/n191 ), 
	.A1(FE_OCPUNCON1077_FE_OFN459_offset_0_), 
	.A0(n2578));
   NAND2BX1TS U1081 (.Y(\add_x_22_3/n24 ), 
	.B(\add_x_22_3/n59 ), 
	.AN(\add_x_22_3/n26 ));
   NAND3X1TS U1082 (.Y(n1288), 
	.C(\add_x_22_5/n77 ), 
	.B(\addr_calc/iir_write_calc/count[14] ), 
	.A(FE_OFN229_addr_calc_iir_write_calc_count_15_));
   NOR3X1TS U1083 (.Y(\add_x_22_5/n59 ), 
	.C(n1288), 
	.B(\add_x_22_5/n69 ), 
	.A(FE_OFN149_add_x_22_5_n94));
   NOR4XLTS U1084 (.Y(n1289), 
	.D(\addr_calc/fft_write_calc/count[16] ), 
	.C(n1976), 
	.B(n1927), 
	.A(\addr_calc/fft_write_calc/count[14] ));
   NOR4X1TS U1085 (.Y(n1290), 
	.D(n1932), 
	.C(\addr_calc/fft_write_calc/count[11] ), 
	.B(\addr_calc/fft_write_calc/count[0] ), 
	.A(n2023));
   NAND4X1TS U1086 (.Y(n1291), 
	.D(n846), 
	.C(n847), 
	.B(n1290), 
	.A(n1289));
   NAND4X2TS U1087 (.Y(n1292), 
	.D(n842), 
	.C(n843), 
	.B(n844), 
	.A(n845));
   NOR2X2TS U1088 (.Y(n2796), 
	.B(n1292), 
	.A(n1291));
   CLKINVX1TS U1089 (.Y(n1293), 
	.A(n1607));
   CLKINVX1TS U1090 (.Y(n1294), 
	.A(FE_OFN144_add_x_19_5_n59));
   AOI32X1TS U1091 (.Y(n1606), 
	.B1(n1294), 
	.B0(n1607), 
	.A2(FE_OFN144_add_x_19_5_n59), 
	.A1(n1293), 
	.A0(\add_x_19_5/n58 ));
   NOR4X1TS U1092 (.Y(n1295), 
	.D(n1972), 
	.C(n2058), 
	.B(\addr_calc/fft_read_calc/count[12] ), 
	.A(n1970));
   NOR4X1TS U1093 (.Y(n1296), 
	.D(n2554), 
	.C(n1967), 
	.B(\addr_calc/fft_read_calc/count[14] ), 
	.A(\addr_calc/fft_read_calc/count[15] ));
   NAND4X1TS U1094 (.Y(n1297), 
	.D(n1296), 
	.C(n1295), 
	.B(n833), 
	.A(n832));
   NAND4X2TS U1095 (.Y(n1298), 
	.D(n831), 
	.C(n830), 
	.B(n829), 
	.A(n828));
   CLKINVX1TS U1099 (.Y(n1301), 
	.A(\add_x_19_3/n129 ));
   OAI2BB1X1TS U1101 (.Y(n1303), 
	.B0(\add_x_19_5/n176 ), 
	.A1N(\add_x_19_5/n219 ), 
	.A0N(n1818));
   CLKINVX1TS U1102 (.Y(n1304), 
	.A(\add_x_19_5/n171 ));
   OAI21XLTS U1103 (.Y(n1305), 
	.B0(n1303), 
	.A1(n1304), 
	.A0(FE_OCPN1225_add_x_19_5_n170));
   OAI31X4TS U1104 (.Y(\addr_calc/iir_write_addr[5] ), 
	.B0(n1305), 
	.A2(n1304), 
	.A1(n1303), 
	.A0(FE_OCPN1225_add_x_19_5_n170));
   OAI2BB1X4TS U1105 (.Y(n1306), 
	.B0(\add_x_19_5/n145 ), 
	.A1N(\add_x_19_5/n213 ), 
	.A0N(\add_x_19_5/n146 ));
   CLKINVX1TS U1106 (.Y(n1307), 
	.A(\add_x_19_5/n140 ));
   OAI21X2TS U1107 (.Y(n1308), 
	.B0(n1306), 
	.A1(n1307), 
	.A0(\add_x_19_5/n139 ));
   OAI31X2TS U1108 (.Y(\addr_calc/iir_write_addr[11] ), 
	.B0(n1308), 
	.A2(n1307), 
	.A1(n1306), 
	.A0(\add_x_19_5/n139 ));
   NAND2BX1TS U1109 (.Y(n1309), 
	.B(\add_x_19_5/n67 ), 
	.AN(\add_x_19_5/n66 ));
   XOR2X4TS U1110 (.Y(\addr_calc/iir_write_addr[24] ), 
	.B(n1309), 
	.A(FE_OCPN1229_add_x_19_5_n68));
   NAND2BX1TS U1111 (.Y(n1310), 
	.B(\add_x_19_0/n166 ), 
	.AN(\add_x_19_0/n165 ));
   XOR2X4TS U1112 (.Y(\addr_calc/fft_read_addr[6] ), 
	.B(n1310), 
	.A(\add_x_19_0/n167 ));
   OAI2BB1X4TS U1113 (.Y(n1311), 
	.B0(\add_x_19_0/n145 ), 
	.A1N(\add_x_19_0/n213 ), 
	.A0N(\add_x_19_0/n146 ));
   CLKINVX1TS U1114 (.Y(n1312), 
	.A(\add_x_19_0/n140 ));
   OAI21X1TS U1117 (.Y(n1314), 
	.B0(\add_x_19_3/n185 ), 
	.A1(\add_x_19_3/n186 ), 
	.A0(\add_x_19_3/n184 ));
   CLKINVX1TS U1118 (.Y(n1315), 
	.A(\add_x_19_3/n182 ));
   OAI21X1TS U1119 (.Y(n1316), 
	.B0(n1314), 
	.A1(n1315), 
	.A0(FE_OCPN1255_add_x_19_3_n181));
   OAI31X2TS U1120 (.Y(\addr_calc/fir_write_addr[3] ), 
	.B0(n1316), 
	.A2(n1315), 
	.A1(n1314), 
	.A0(FE_OCPN1255_add_x_19_3_n181));
   OA21XLTS U1121 (.Y(\addr_calc/iir_read_addr[0] ), 
	.B0(\add_x_19_4/n191 ), 
	.A1(FE_OCPUNCON1077_FE_OFN459_offset_0_), 
	.A0(n2580));
   NOR4XLTS U1122 (.Y(n1317), 
	.D(instruction[15]), 
	.C(instruction[13]), 
	.B(instruction[10]), 
	.A(instruction[14]));
   NOR4XLTS U1123 (.Y(n1318), 
	.D(instruction[21]), 
	.C(instruction[22]), 
	.B(instruction[20]), 
	.A(instruction[24]));
   NOR4BBX1TS U1124 (.Y(n1319), 
	.D(instruction[16]), 
	.C(instruction[17]), 
	.BN(n2093), 
	.AN(n2108));
   NAND4X1TS U1125 (.Y(n908), 
	.D(n1319), 
	.C(n1318), 
	.B(n802), 
	.A(n1317));
   NAND4BX1TS U1126 (.Y(\add_x_22_5/n94 ), 
	.D(\addr_calc/iir_write_calc/count[6] ), 
	.C(n1683), 
	.B(\add_x_22_5/n111 ), 
	.AN(\add_x_22_5/n103 ));
   NAND4BX2TS U1127 (.Y(\add_x_22_3/n94 ), 
	.D(FE_OFN254_addr_calc_fir_write_calc_count_6_), 
	.C(n1869), 
	.B(\add_x_22_3/n111 ), 
	.AN(\add_x_22_3/n103 ));
   NAND2BX1TS U1128 (.Y(\add_x_22_2/n24 ), 
	.B(FE_OFN147_add_x_22_2_n59), 
	.AN(\add_x_22_2/n26 ));
   NAND2BX1TS U1129 (.Y(\add_x_22_4/n85 ), 
	.B(\add_x_22_4/n93 ), 
	.AN(\add_x_22_4/n87 ));
   NAND2BX1TS U1132 (.Y(n1321), 
	.B(\add_x_19_1/n59 ), 
	.AN(\add_x_19_1/n58 ));
   NAND2BX1TS U1133 (.Y(n1322), 
	.B(\add_x_19_1/n101 ), 
	.AN(\add_x_19_1/n100 ));
   XOR2X4TS U1134 (.Y(\addr_calc/fft_write_addr[18] ), 
	.B(n1322), 
	.A(\add_x_19_1/n102 ));
   NAND2BX1TS U1135 (.Y(n1323), 
	.B(\add_x_19_5/n82 ), 
	.AN(\add_x_19_5/n81 ));
   XNOR2X1TS U1137 (.Y(n1324), 
	.B(\add_x_22_1/n118 ), 
	.A(\add_x_22_1/n117 ));
   AO22X4TS U1138 (.Y(n1064), 
	.B1(n1324), 
	.B0(FE_OFN34_n2795), 
	.A1(n2032), 
	.A0(FE_OFN25_n2797));
   NAND2BXLTS U1139 (.Y(n1325), 
	.B(FE_OFN142_add_x_19_2_n59), 
	.AN(\add_x_19_2/n58 ));
   NAND2BX1TS U1140 (.Y(n1326), 
	.B(\add_x_19_5/n155 ), 
	.AN(\add_x_19_5/n154 ));
   XOR2X1TS U1141 (.Y(\addr_calc/iir_write_addr[8] ), 
	.B(n1326), 
	.A(\add_x_19_5/n156 ));
   NAND2BX1TS U1142 (.Y(n1327), 
	.B(\add_x_19_5/n132 ), 
	.AN(\add_x_19_5/n131 ));
   XOR2X2TS U1143 (.Y(\addr_calc/iir_write_addr[12] ), 
	.B(n1327), 
	.A(\add_x_19_5/n133 ));
   OAI2BB1X4TS U1144 (.Y(n1328), 
	.B0(\add_x_19_3/n145 ), 
	.A1N(\add_x_19_3/n213 ), 
	.A0N(\add_x_19_3/n146 ));
   CLKINVX1TS U1145 (.Y(n1329), 
	.A(\add_x_19_3/n140 ));
   OAI21X1TS U1146 (.Y(n1330), 
	.B0(n1328), 
	.A1(n1329), 
	.A0(FE_OCPN1906_add_x_19_3_n139));
   OAI31X2TS U1147 (.Y(\addr_calc/fir_write_addr[11] ), 
	.B0(n1330), 
	.A2(n1329), 
	.A1(n1328), 
	.A0(FE_OCPN1906_add_x_19_3_n139));
   CLKINVX1TS U1149 (.Y(n1332), 
	.A(\add_x_19_3/n106 ));
   OAI21X1TS U1150 (.Y(n1333), 
	.B0(n1331), 
	.A1(n1332), 
	.A0(\add_x_19_3/n105 ));
   OAI31X2TS U1151 (.Y(\addr_calc/fir_write_addr[17] ), 
	.B0(n1333), 
	.A2(n1332), 
	.A1(n1331), 
	.A0(\add_x_19_3/n105 ));
   NAND2BXLTS U1152 (.Y(n1334), 
	.B(\add_x_19_3/n67 ), 
	.AN(\add_x_19_3/n66 ));
   OAI2BB1X1TS U1154 (.Y(n1335), 
	.B0(\add_x_19_2/n176 ), 
	.A1N(\add_x_19_2/n219 ), 
	.A0N(\add_x_19_2/n177 ));
   CLKINVX1TS U1155 (.Y(n1336), 
	.A(\add_x_19_2/n171 ));
   OAI21XLTS U1156 (.Y(n1337), 
	.B0(n1335), 
	.A1(n1336), 
	.A0(\add_x_19_2/n170 ));
   OAI31XLTS U1157 (.Y(\addr_calc/fir_read_addr[5] ), 
	.B0(n1337), 
	.A2(n1336), 
	.A1(n1335), 
	.A0(\add_x_19_2/n170 ));
   OAI21X1TS U1158 (.Y(n1338), 
	.B0(\add_x_19_4/n166 ), 
	.A1(\add_x_19_4/n167 ), 
	.A0(\add_x_19_4/n165 ));
   CLKINVX1TS U1159 (.Y(n1339), 
	.A(\add_x_19_4/n163 ));
   OAI21X2TS U1160 (.Y(n1340), 
	.B0(n1338), 
	.A1(n1339), 
	.A0(FE_OCPN1221_add_x_19_4_n162));
   OAI31X2TS U1161 (.Y(\addr_calc/iir_read_addr[7] ), 
	.B0(n1340), 
	.A2(n1339), 
	.A1(n1338), 
	.A0(FE_OCPN1221_add_x_19_4_n162));
   OAI21X1TS U1162 (.Y(n1341), 
	.B0(\add_x_19_2/n155 ), 
	.A1(\add_x_19_2/n156 ), 
	.A0(\add_x_19_2/n154 ));
   INVXLTS U1163 (.Y(n1342), 
	.A(\add_x_19_2/n152 ));
   OAI21XLTS U1164 (.Y(n1343), 
	.B0(n1341), 
	.A1(n1342), 
	.A0(\add_x_19_2/n151 ));
   OAI31X1TS U1165 (.Y(\addr_calc/fir_read_addr[9] ), 
	.B0(n1343), 
	.A2(n1342), 
	.A1(n1341), 
	.A0(\add_x_19_2/n151 ));
   NAND2BX1TS U1166 (.Y(n1344), 
	.B(\add_x_19_5/n185 ), 
	.AN(\add_x_19_5/n184 ));
   XOR2X1TS U1167 (.Y(\addr_calc/iir_write_addr[2] ), 
	.B(n1344), 
	.A(\add_x_19_5/n186 ));
   NAND2BX1TS U1168 (.Y(n1345), 
	.B(\add_x_19_2/n189 ), 
	.AN(\add_x_19_2/n188 ));
   XOR2X1TS U1169 (.Y(\addr_calc/fir_read_addr[1] ), 
	.B(n1345), 
	.A(\add_x_19_2/n191 ));
   OAI21X1TS U1170 (.Y(n1346), 
	.B0(\add_x_19_2/n185 ), 
	.A1(\add_x_19_2/n186 ), 
	.A0(\add_x_19_2/n184 ));
   CLKINVX1TS U1171 (.Y(n1347), 
	.A(\add_x_19_2/n182 ));
   OAI21X1TS U1172 (.Y(n1348), 
	.B0(n1346), 
	.A1(n1347), 
	.A0(FE_OCPN1220_add_x_19_2_n181));
   OAI31X1TS U1173 (.Y(\addr_calc/fir_read_addr[3] ), 
	.B0(n1348), 
	.A2(n1347), 
	.A1(n1346), 
	.A0(FE_OCPN1220_add_x_19_2_n181));
   OA21XLTS U1174 (.Y(\addr_calc/fir_write_addr[0] ), 
	.B0(\add_x_19_3/n191 ), 
	.A1(FE_OFN461_offset_0_), 
	.A0(FE_OFN252_addr_calc_fir_write_calc_count_0_));
   NAND4BX1TS U1175 (.Y(n1349), 
	.D(\add_x_22_1/n77 ), 
	.C(\addr_calc/fft_write_calc/count[15] ), 
	.B(FE_OFN259_addr_calc_fft_write_calc_count_14_), 
	.AN(\add_x_22_1/n69 ));
   NOR2X2TS U1176 (.Y(\add_x_22_1/n59 ), 
	.B(n1349), 
	.A(\add_x_22_1/n94 ));
   NAND2BX1TS U1177 (.Y(\add_x_22_5/n24 ), 
	.B(FE_OFN148_add_x_22_5_n59), 
	.AN(\add_x_22_5/n26 ));
   NAND4BX2TS U1178 (.Y(\add_x_22_4/n94 ), 
	.D(\addr_calc/iir_read_calc/count[6] ), 
	.C(FE_OFN246_addr_calc_iir_read_calc_count_7_), 
	.B(\add_x_22_4/n111 ), 
	.AN(\add_x_22_4/n103 ));
   NAND2BX1TS U1179 (.Y(\add_x_22_0/n85 ), 
	.B(\add_x_22_0/n93 ), 
	.AN(\add_x_22_0/n87 ));
   AND4X1TS U1180 (.Y(n1350), 
	.D(instruction[30]), 
	.C(instruction[29]), 
	.B(instruction[28]), 
	.A(instruction[26]));
   AND3X1TS U1181 (.Y(n802), 
	.C(n1350), 
	.B(instruction[27]), 
	.A(instruction[31]));
   NAND2BX1TS U1182 (.Y(n1351), 
	.B(\add_x_19_0/n101 ), 
	.AN(\add_x_19_0/n100 ));
   NAND2BX1TS U1184 (.Y(n1352), 
	.B(\add_x_19_2/n82 ), 
	.AN(\add_x_19_2/n81 ));
   XOR2X4TS U1185 (.Y(\addr_calc/fir_read_addr[22] ), 
	.B(n1352), 
	.A(FE_OCPN1362_add_x_19_2_n83));
   XNOR2X1TS U1186 (.Y(n1353), 
	.B(\add_x_22_1/n121 ), 
	.A(FE_OFN260_addr_calc_fft_write_calc_count_0_));
   AO22X4TS U1187 (.Y(n1065), 
	.B1(n1353), 
	.B0(FE_OFN34_n2795), 
	.A1(n1941), 
	.A0(FE_OFN25_n2797));
   NAND2BX1TS U1188 (.Y(n1354), 
	.B(FE_OFN144_add_x_19_5_n59), 
	.AN(\add_x_19_5/n58 ));
   CLKXOR2X4TS U1189 (.Y(\addr_calc/iir_write_addr[26] ), 
	.B(n1354), 
	.A(\add_x_19_5/n60 ));
   NAND2BX1TS U1190 (.Y(n1355), 
	.B(\add_x_19_4/n59 ), 
	.AN(\add_x_19_4/n58 ));
   XOR2X4TS U1191 (.Y(\addr_calc/iir_read_addr[26] ), 
	.B(n1355), 
	.A(\add_x_19_4/n60 ));
   OAI2BB1X1TS U1193 (.Y(n1357), 
	.B0(n1586), 
	.A1N(FE_OFN340_offset_31_), 
	.A0N(FE_OFN234_addr_calc_iir_read_calc_count_31_));
   AOI21X4TS U1194 (.Y(n1358), 
	.B0(n1589), 
	.A1(n2629), 
	.A0(FE_OFN531_add_x_19_5_n43));
   NAND2XLTS U1195 (.Y(n1359), 
	.B(\add_x_19_5/n37 ), 
	.A(n1533));
   NAND2BX1TS U1197 (.Y(n1360), 
	.B(\add_x_19_5/n124 ), 
	.AN(\add_x_19_5/n123 ));
   NAND2BX1TS U1199 (.Y(n1361), 
	.B(\add_x_19_5/n90 ), 
	.AN(\add_x_19_5/n89 ));
   XOR2X4TS U1200 (.Y(\addr_calc/iir_write_addr[20] ), 
	.B(n1361), 
	.A(\add_x_19_5/n91 ));
   NAND2BX1TS U1201 (.Y(n1362), 
	.B(\add_x_19_4/n155 ), 
	.AN(\add_x_19_4/n154 ));
   CLKXOR2X2TS U1202 (.Y(\addr_calc/iir_read_addr[8] ), 
	.B(n1362), 
	.A(FE_OCP_RBN1925_add_x_19_4_n157));
   NAND2BX1TS U1203 (.Y(n1363), 
	.B(\add_x_19_2/n132 ), 
	.AN(\add_x_19_2/n131 ));
   NAND2BXLTS U1205 (.Y(n1364), 
	.B(\add_x_19_2/n67 ), 
	.AN(\add_x_19_2/n66 ));
   XOR2X4TS U1206 (.Y(\addr_calc/fir_read_addr[24] ), 
	.B(n1364), 
	.A(\add_x_19_2/n68 ));
   NAND2BX1TS U1207 (.Y(n1365), 
	.B(\add_x_19_0/n185 ), 
	.AN(\add_x_19_0/n184 ));
   XOR2X1TS U1208 (.Y(\addr_calc/fft_read_addr[2] ), 
	.B(n1365), 
	.A(\add_x_19_0/n186 ));
   CLKINVX1TS U1209 (.Y(n1366), 
	.A(\add_x_19_0/n171 ));
   OAI2BB1X1TS U1210 (.Y(n1367), 
	.B0(\add_x_19_0/n176 ), 
	.A1N(\add_x_19_0/n219 ), 
	.A0N(\add_x_19_0/n177 ));
   OAI21XLTS U1211 (.Y(n1368), 
	.B0(n1367), 
	.A1(n1366), 
	.A0(\add_x_19_0/n170 ));
   OAI31X4TS U1212 (.Y(\addr_calc/fft_read_addr[5] ), 
	.B0(n1368), 
	.A2(n1366), 
	.A1(n1367), 
	.A0(\add_x_19_0/n170 ));
   OAI21X1TS U1213 (.Y(n1369), 
	.B0(\add_x_19_5/n166 ), 
	.A1(\add_x_19_5/n167 ), 
	.A0(\add_x_19_5/n165 ));
   CLKINVX1TS U1214 (.Y(n1370), 
	.A(\add_x_19_5/n163 ));
   OAI21X1TS U1215 (.Y(n1371), 
	.B0(n1369), 
	.A1(n1370), 
	.A0(FE_OCPN1222_add_x_19_5_n162));
   OAI31X1TS U1216 (.Y(\addr_calc/iir_write_addr[7] ), 
	.B0(n1371), 
	.A2(n1370), 
	.A1(n1369), 
	.A0(FE_OCPN1222_add_x_19_5_n162));
   NAND2X1TS U1217 (.Y(n1372), 
	.B(\add_x_19_3/n111 ), 
	.A(\add_x_19_3/n207 ));
   XNOR2X1TS U1218 (.Y(\addr_calc/fir_write_addr[16] ), 
	.B(FE_OCP_RBN1378_add_x_19_3_n113), 
	.A(n1372));
   OAI21X2TS U1219 (.Y(n1373), 
	.B0(\add_x_19_1/n166 ), 
	.A1(\add_x_19_1/n167 ), 
	.A0(\add_x_19_1/n165 ));
   CLKINVX1TS U1220 (.Y(n1374), 
	.A(\add_x_19_1/n163 ));
   OAI21X1TS U1221 (.Y(n1375), 
	.B0(n1373), 
	.A1(n1374), 
	.A0(\add_x_19_1/n162 ));
   OAI31X4TS U1222 (.Y(\addr_calc/fft_write_addr[7] ), 
	.B0(n1375), 
	.A2(n1374), 
	.A1(n1373), 
	.A0(\add_x_19_1/n162 ));
   OAI21X1TS U1223 (.Y(n1376), 
	.B0(\add_x_19_1/n155 ), 
	.A1(FE_OCP_RBN1956_FE_OFN520_add_x_19_1_n157), 
	.A0(\add_x_19_1/n154 ));
   CLKINVX1TS U1224 (.Y(n1377), 
	.A(\add_x_19_1/n152 ));
   OAI21XLTS U1225 (.Y(n1378), 
	.B0(n1376), 
	.A1(n1377), 
	.A0(\add_x_19_1/n151 ));
   OAI31X4TS U1226 (.Y(\addr_calc/fft_write_addr[9] ), 
	.B0(n1378), 
	.A2(n1377), 
	.A1(n1376), 
	.A0(\add_x_19_1/n151 ));
   NAND2BX1TS U1227 (.Y(n1379), 
	.B(\add_x_19_3/n189 ), 
	.AN(\add_x_19_3/n188 ));
   XOR2X1TS U1228 (.Y(\addr_calc/fir_write_addr[1] ), 
	.B(n1379), 
	.A(\add_x_19_3/n191 ));
   OAI21X1TS U1229 (.Y(n1380), 
	.B0(\add_x_19_1/n185 ), 
	.A1(FE_OCP_RBN1955_add_x_19_1_n187), 
	.A0(\add_x_19_1/n184 ));
   CLKINVX1TS U1230 (.Y(n1381), 
	.A(\add_x_19_1/n182 ));
   OAI21XLTS U1231 (.Y(n1382), 
	.B0(n1380), 
	.A1(n1381), 
	.A0(FE_OCPN1223_add_x_19_1_n181));
   OAI31X1TS U1232 (.Y(\addr_calc/fft_write_addr[3] ), 
	.B0(n1382), 
	.A2(n1381), 
	.A1(n1380), 
	.A0(FE_OCPN1223_add_x_19_1_n181));
   OA21XLTS U1233 (.Y(\addr_calc/fir_read_addr[0] ), 
	.B0(\add_x_19_2/n191 ), 
	.A1(FE_OCPUNCON1068_offset_0_), 
	.A0(n2007));
   NAND4BX1TS U1234 (.Y(\add_x_22_2/n26 ), 
	.D(\add_x_22_2/n43 ), 
	.C(n1691), 
	.B(n2558), 
	.AN(\add_x_22_2/n35 ));
   NAND4BX1TS U1235 (.Y(\add_x_22_0/n26 ), 
	.D(\add_x_22_0/n43 ), 
	.C(\addr_calc/fft_read_calc/count[22] ), 
	.B(\addr_calc/fft_read_calc/count[23] ), 
	.AN(\add_x_22_0/n35 ));
   NAND2BX1TS U1236 (.Y(\add_x_22_4/n24 ), 
	.B(FE_OFN150_add_x_22_4_n59), 
	.AN(\add_x_22_4/n26 ));
   NAND2BX1TS U1237 (.Y(\add_x_22_1/n24 ), 
	.B(\add_x_22_1/n59 ), 
	.AN(\add_x_22_1/n26 ));
   NAND2BX1TS U1238 (.Y(\add_x_22_3/n85 ), 
	.B(\add_x_22_3/n93 ), 
	.AN(\add_x_22_3/n87 ));
   NAND2BX1TS U1239 (.Y(\add_x_22_2/n85 ), 
	.B(\add_x_22_2/n93 ), 
	.AN(\add_x_22_2/n87 ));
   NAND2BX1TS U1240 (.Y(n884), 
	.B(n902), 
	.AN(n2311));
   XOR2X1TS U1241 (.Y(n1383), 
	.B(n2031), 
	.A(\add_x_22_4/n34 ));
   AO22X1TS U1242 (.Y(n949), 
	.B1(FE_OFN91_n1192), 
	.B0(n2031), 
	.A1(n1383), 
	.A0(FE_OFN79_n2787));
   NAND2BX2TS U1244 (.Y(n1385), 
	.B(\add_x_19_1/n106 ), 
	.AN(\add_x_19_1/n105 ));
   NAND2BX1TS U1246 (.Y(n1386), 
	.B(\add_x_19_1/n124 ), 
	.AN(\add_x_19_1/n123 ));
   XOR2X2TS U1247 (.Y(\addr_calc/fft_write_addr[14] ), 
	.B(n1386), 
	.A(\add_x_19_1/n125 ));
   NAND2BXLTS U1248 (.Y(n1387), 
	.B(\add_x_19_5/n101 ), 
	.AN(\add_x_19_5/n100 ));
   NAND2BX1TS U1250 (.Y(n1388), 
	.B(\add_x_19_4/n101 ), 
	.AN(\add_x_19_4/n100 ));
   NOR2X1TS U1252 (.Y(n1389), 
	.B(\add_x_22_1/n85 ), 
	.A(\add_x_22_1/n84 ));
   XNOR2X1TS U1253 (.Y(n1390), 
	.B(n1930), 
	.A(n1389));
   AO22X1TS U1254 (.Y(n1055), 
	.B1(n1390), 
	.B0(n2795), 
	.A1(n1667), 
	.A0(FE_OCPN1911_FE_OFN17_n2797));
   NAND2BXLTS U1255 (.Y(n1391), 
	.B(\add_x_19_3/n82 ), 
	.AN(\add_x_19_3/n81 ));
   NAND2BX1TS U1257 (.Y(n1392), 
	.B(\add_x_19_0/n59 ), 
	.AN(\add_x_19_0/n58 ));
   XOR2X4TS U1258 (.Y(\addr_calc/fft_read_addr[26] ), 
	.B(n1392), 
	.A(\add_x_19_0/n60 ));
   NAND2BX2TS U1259 (.Y(n1393), 
	.B(\add_x_19_0/n90 ), 
	.AN(\add_x_19_0/n89 ));
   OAI2BB2XLTS U1260 (.Y(n1034), 
	.B1(n1394), 
	.B0(n2794), 
	.A1N(n2794), 
	.A0N(FE_OFN517_addr_calc_fft_read_calc_count_0_));
   NAND2X1TS U1261 (.Y(n1395), 
	.B(FE_OFN282_addr_calc_fir_write_calc_count_20_), 
	.A(\add_x_22_3/n41 ));
   XOR2X1TS U1262 (.Y(n1396), 
	.B(n1395), 
	.A(n1891));
   AO22X1TS U1263 (.Y(n1109), 
	.B1(n1396), 
	.B0(n1762), 
	.A1(FE_OCPUNCON1087_n2805), 
	.A0(\addr_calc/fir_write_calc/count[21] ));
   CLKINVX1TS U1265 (.Y(n1398), 
	.A(\add_x_19_4/n171 ));
   OAI31X4TS U1267 (.Y(\addr_calc/iir_read_addr[5] ), 
	.B0(n1399), 
	.A2(n1398), 
	.A1(n1397), 
	.A0(\add_x_19_4/n170 ));
   NAND2BX1TS U1268 (.Y(n1400), 
	.B(\add_x_19_4/n124 ), 
	.AN(\add_x_19_4/n123 ));
   XOR2X4TS U1269 (.Y(\addr_calc/iir_read_addr[14] ), 
	.B(n1400), 
	.A(\add_x_19_4/n125 ));
   NAND2BX1TS U1270 (.Y(n1401), 
	.B(\add_x_19_3/n132 ), 
	.AN(\add_x_19_3/n131 ));
   CLKXOR2X2TS U1271 (.Y(\addr_calc/fir_write_addr[12] ), 
	.B(n1401), 
	.A(\add_x_19_3/n133 ));
   AOI21X2TS U1272 (.Y(n1402), 
	.B0(\add_x_19_2/n143 ), 
	.A1(\add_x_19_2/n213 ), 
	.A0(\add_x_19_2/n146 ));
   NAND2X1TS U1273 (.Y(n1403), 
	.B(\add_x_19_2/n140 ), 
	.A(\add_x_19_2/n212 ));
   XOR2X4TS U1274 (.Y(\addr_calc/fir_read_addr[11] ), 
	.B(n1403), 
	.A(n1402));
   NAND2BX4TS U1275 (.Y(n1404), 
	.B(\add_x_19_2/n90 ), 
	.AN(\add_x_19_2/n89 ));
   NAND2BX1TS U1276 (.Y(n1405), 
	.B(\add_x_19_1/n155 ), 
	.AN(\add_x_19_1/n154 ));
   NAND2BX1TS U1277 (.Y(n1406), 
	.B(\add_x_19_1/n67 ), 
	.AN(\add_x_19_1/n66 ));
   NAND2BX4TS U1278 (.Y(n1407), 
	.B(\add_x_19_0/n132 ), 
	.AN(\add_x_19_0/n131 ));
   XOR2X4TS U1279 (.Y(\addr_calc/fft_read_addr[12] ), 
	.B(n1407), 
	.A(\add_x_19_0/n133 ));
   NAND2X1TS U1280 (.Y(n1408), 
	.B(\add_x_19_5/n42 ), 
	.A(n2629));
   OAI21X1TS U1282 (.Y(n1409), 
	.B0(\add_x_19_4/n155 ), 
	.A1(\add_x_19_4/n154 ), 
	.A0(FE_OCP_RBN1925_add_x_19_4_n157));
   CLKINVX1TS U1283 (.Y(n1410), 
	.A(\add_x_19_4/n152 ));
   OAI21X1TS U1286 (.Y(n1412), 
	.B0(\add_x_19_3/n166 ), 
	.A1(\add_x_19_3/n167 ), 
	.A0(\add_x_19_3/n165 ));
   OAI21X1TS U1288 (.Y(n1414), 
	.B0(n1412), 
	.A1(FE_OCP_RBN1788_add_x_19_3_n163), 
	.A0(FE_OCPN1256_add_x_19_3_n162));
   OAI31X1TS U1289 (.Y(\addr_calc/fir_write_addr[7] ), 
	.B0(n1414), 
	.A2(FE_OCP_RBN1788_add_x_19_3_n163), 
	.A1(n1412), 
	.A0(FE_OCPN1256_add_x_19_3_n162));
   NAND2X1TS U1290 (.Y(n1415), 
	.B(\add_x_19_3/n42 ), 
	.A(n2631));
   XNOR2X4TS U1291 (.Y(\addr_calc/fir_write_addr[29] ), 
	.B(\add_x_19_3/n43 ), 
	.A(n1415));
   NAND2X2TS U1292 (.Y(n1416), 
	.B(\add_x_19_2/n111 ), 
	.A(\add_x_19_2/n207 ));
   OAI21X1TS U1294 (.Y(n1417), 
	.B0(\add_x_19_0/n155 ), 
	.A1(\add_x_19_0/n156 ), 
	.A0(\add_x_19_0/n154 ));
   CLKINVX1TS U1295 (.Y(n1418), 
	.A(\add_x_19_0/n152 ));
   OAI21X1TS U1296 (.Y(n1419), 
	.B0(n1417), 
	.A1(n1418), 
	.A0(\add_x_19_0/n151 ));
   NAND2X1TS U1298 (.Y(n1420), 
	.B(\add_x_19_0/n111 ), 
	.A(\add_x_19_0/n207 ));
   NAND2BX1TS U1300 (.Y(n1421), 
	.B(\add_x_19_2/n185 ), 
	.AN(\add_x_19_2/n184 ));
   XOR2X1TS U1301 (.Y(\addr_calc/fir_read_addr[2] ), 
	.B(n1421), 
	.A(\add_x_19_2/n186 ));
   NAND2BX1TS U1302 (.Y(n1422), 
	.B(\add_x_19_0/n189 ), 
	.AN(\add_x_19_0/n188 ));
   XOR2X1TS U1303 (.Y(\addr_calc/fft_read_addr[1] ), 
	.B(n1422), 
	.A(\add_x_19_0/n191 ));
   CLKINVX1TS U1304 (.Y(n1423), 
	.A(\add_x_19_0/n182 ));
   OAI21X1TS U1305 (.Y(n1424), 
	.B0(\add_x_19_0/n185 ), 
	.A1(\add_x_19_0/n186 ), 
	.A0(\add_x_19_0/n184 ));
   OAI21XLTS U1306 (.Y(n1425), 
	.B0(n1424), 
	.A1(n1423), 
	.A0(FE_OCPN1189_add_x_19_0_n181));
   OAI31X1TS U1307 (.Y(\addr_calc/fft_read_addr[3] ), 
	.B0(n1425), 
	.A2(n1423), 
	.A1(n1424), 
	.A0(FE_OCPN1189_add_x_19_0_n181));
   OA21XLTS U1308 (.Y(\addr_calc/fft_write_addr[0] ), 
	.B0(\add_x_19_1/n191 ), 
	.A1(FE_OFN459_offset_0_), 
	.A0(FE_OFN260_addr_calc_fft_write_calc_count_0_));
   NAND4BX1TS U1309 (.Y(\add_x_22_5/n26 ), 
	.D(\add_x_22_5/n43 ), 
	.C(n2579), 
	.B(\addr_calc/iir_write_calc/count[23] ), 
	.AN(\add_x_22_5/n35 ));
   NAND2BX1TS U1310 (.Y(\add_x_22_0/n24 ), 
	.B(\add_x_22_0/n59 ), 
	.AN(\add_x_22_0/n26 ));
   NAND3BX2TS U1311 (.Y(\DP_OP_158_296_6262/n1834 ), 
	.C(\DP_OP_158_296_6262/n1837 ), 
	.B(FE_OFN113_DP_OP_158_296_6262_n1791), 
	.AN(\DP_OP_158_296_6262/n1792 ));
   OAI21X2TS U1312 (.Y(n1426), 
	.B0(\add_x_19_5/n56 ), 
	.A1(\add_x_19_5/n59 ), 
	.A0(\add_x_19_5/n55 ));
   AOI21X2TS U1313 (.Y(\add_x_19_5/n52 ), 
	.B0(n1426), 
	.A1(\add_x_19_5/n62 ), 
	.A0(\add_x_19_5/n53 ));
   NAND2BX1TS U1314 (.Y(\add_x_22_5/n85 ), 
	.B(\add_x_22_5/n93 ), 
	.AN(\add_x_22_5/n87 ));
   NAND2BX1TS U1315 (.Y(\add_x_22_1/n85 ), 
	.B(\add_x_22_1/n93 ), 
	.AN(\add_x_22_1/n87 ));
   NAND4BX1TS U1316 (.Y(n1427), 
	.D(\add_x_22_3/n9 ), 
	.C(n1896), 
	.B(\add_x_22_3/n59 ), 
	.AN(\add_x_22_3/n26 ));
   NOR2BX1TS U1317 (.Y(\add_x_22_3/n2 ), 
	.B(n1427), 
	.AN(\addr_calc/fir_write_calc/count[29] ));
   XNOR2X1TS U1318 (.Y(\addr_calc/fir_write_calc/counter/N72 ), 
	.B(n1427), 
	.A(\addr_calc/fir_write_calc/count[29] ));
   NAND4BX1TS U1319 (.Y(n1428), 
	.D(\add_x_22_4/n9 ), 
	.C(n2561), 
	.B(FE_OFN150_add_x_22_4_n59), 
	.AN(\add_x_22_4/n26 ));
   NOR2BX1TS U1320 (.Y(\add_x_22_4/n2 ), 
	.B(n1428), 
	.AN(\addr_calc/iir_read_calc/count[29] ));
   XNOR2X1TS U1321 (.Y(\addr_calc/iir_read_calc/counter/N72 ), 
	.B(n1428), 
	.A(\addr_calc/iir_read_calc/count[29] ));
   NAND4BX1TS U1322 (.Y(n1429), 
	.D(\add_x_22_2/n9 ), 
	.C(\addr_calc/fir_read_calc/count[28] ), 
	.B(FE_OFN147_add_x_22_2_n59), 
	.AN(\add_x_22_2/n26 ));
   NOR2BX1TS U1323 (.Y(\add_x_22_2/n2 ), 
	.B(n1429), 
	.AN(\addr_calc/fir_read_calc/count[29] ));
   XNOR2X1TS U1324 (.Y(\addr_calc/fir_read_calc/counter/N72 ), 
	.B(n1429), 
	.A(\addr_calc/fir_read_calc/count[29] ));
   NAND2BX1TS U1325 (.Y(n1430), 
	.B(\add_x_19_1/n37 ), 
	.AN(\add_x_19_1/n36 ));
   XOR2X2TS U1326 (.Y(\addr_calc/fft_write_addr[30] ), 
	.B(n1430), 
	.A(\add_x_19_1/n38 ));
   NAND2BX2TS U1327 (.Y(n1431), 
	.B(\add_x_19_3/n101 ), 
	.AN(\add_x_19_3/n100 ));
   NAND2BX1TS U1329 (.Y(n1432), 
	.B(\add_x_19_2/n101 ), 
	.AN(\add_x_19_2/n100 ));
   NAND2BX1TS U1331 (.Y(n1433), 
	.B(\add_x_19_4/n82 ), 
	.AN(\add_x_19_4/n81 ));
   NAND2BX1TS U1332 (.Y(n1434), 
	.B(\add_x_19_0/n82 ), 
	.AN(\add_x_19_0/n81 ));
   NAND2BX1TS U1334 (.Y(n1435), 
	.B(FE_OFN143_add_x_19_3_n59), 
	.AN(\add_x_19_3/n58 ));
   XOR2X2TS U1335 (.Y(\addr_calc/fir_write_addr[26] ), 
	.B(n1435), 
	.A(\add_x_19_3/n60 ));
   NAND2BX1TS U1336 (.Y(n1436), 
	.B(\add_x_19_5/n166 ), 
	.AN(\add_x_19_5/n165 ));
   XOR2X1TS U1337 (.Y(\addr_calc/iir_write_addr[6] ), 
	.B(n1436), 
	.A(\add_x_19_5/n167 ));
   NAND2BX1TS U1338 (.Y(n1437), 
	.B(\add_x_19_4/n132 ), 
	.AN(\add_x_19_4/n131 ));
   XOR2X4TS U1339 (.Y(\addr_calc/iir_read_addr[12] ), 
	.B(n1437), 
	.A(\add_x_19_4/n133 ));
   NAND2BXLTS U1340 (.Y(n1438), 
	.B(\add_x_19_3/n90 ), 
	.AN(\add_x_19_3/n89 ));
   NAND2BX1TS U1342 (.Y(n1439), 
	.B(\add_x_19_2/n124 ), 
	.AN(\add_x_19_2/n123 ));
   XOR2X4TS U1343 (.Y(\addr_calc/fir_read_addr[14] ), 
	.B(n1439), 
	.A(\add_x_19_2/n125 ));
   NAND2BX1TS U1344 (.Y(n1440), 
	.B(\add_x_19_1/n132 ), 
	.AN(\add_x_19_1/n131 ));
   XOR2X4TS U1345 (.Y(\addr_calc/fft_write_addr[12] ), 
	.B(n1440), 
	.A(\add_x_19_1/n133 ));
   NAND2BX1TS U1346 (.Y(n1441), 
	.B(\add_x_19_1/n90 ), 
	.AN(\add_x_19_1/n89 ));
   NAND2BX1TS U1347 (.Y(n1442), 
	.B(\add_x_19_0/n124 ), 
	.AN(\add_x_19_0/n123 ));
   CLKXOR2X2TS U1348 (.Y(\addr_calc/fft_read_addr[14] ), 
	.B(n1442), 
	.A(\add_x_19_0/n125 ));
   NAND2X1TS U1349 (.Y(n1443), 
	.B(\add_x_19_4/n111 ), 
	.A(\add_x_19_4/n207 ));
   XNOR2X2TS U1350 (.Y(\addr_calc/iir_read_addr[16] ), 
	.B(n1443), 
	.A(FE_OCPN1226_add_x_19_4_n112));
   NAND2X1TS U1351 (.Y(n1444), 
	.B(\add_x_19_2/n145 ), 
	.A(\add_x_19_2/n213 ));
   XNOR2X1TS U1352 (.Y(\addr_calc/fir_read_addr[10] ), 
	.B(\add_x_19_2/n146 ), 
	.A(n1444));
   NAND2X1TS U1353 (.Y(n1445), 
	.B(\add_x_19_2/n42 ), 
	.A(n2633));
   XNOR2X4TS U1354 (.Y(\addr_calc/fir_read_addr[29] ), 
	.B(\add_x_19_2/n43 ), 
	.A(n1445));
   NAND2X1TS U1355 (.Y(n1446), 
	.B(\add_x_19_1/n145 ), 
	.A(\add_x_19_1/n213 ));
   NAND2X2TS U1356 (.Y(n1447), 
	.B(\add_x_19_1/n111 ), 
	.A(\add_x_19_1/n207 ));
   OAI21X1TS U1357 (.Y(n1448), 
	.B0(\add_x_19_0/n166 ), 
	.A1(\add_x_19_0/n167 ), 
	.A0(\add_x_19_0/n165 ));
   CLKINVX1TS U1358 (.Y(n1449), 
	.A(\add_x_19_0/n163 ));
   OAI21X1TS U1359 (.Y(n1450), 
	.B0(n1448), 
	.A1(n1449), 
	.A0(FE_OCPN1257_add_x_19_0_n162));
   OAI31X1TS U1360 (.Y(\addr_calc/fft_read_addr[7] ), 
	.B0(n1450), 
	.A2(n1449), 
	.A1(n1448), 
	.A0(FE_OCPN1257_add_x_19_0_n162));
   NAND2X1TS U1361 (.Y(n1451), 
	.B(\add_x_19_0/n42 ), 
	.A(n2628));
   NAND3X1TS U1363 (.Y(n1452), 
	.C(n801), 
	.B(FE_OFN336_instruction_0_), 
	.A(n802));
   AOI211X1TS U1364 (.Y(\pla_top/N59 ), 
	.C0(n1452), 
	.B0(acc_done), 
	.A1(n2311), 
	.A0(FE_OFN335_instruction_2_));
   NAND2BX1TS U1365 (.Y(n1453), 
	.B(\add_x_19_1/n189 ), 
	.AN(\add_x_19_1/n188 ));
   XOR2X1TS U1366 (.Y(\addr_calc/fft_write_addr[1] ), 
	.B(n1453), 
	.A(\add_x_19_1/n191 ));
   NAND2BX1TS U1367 (.Y(n1454), 
	.B(\add_x_19_1/n185 ), 
	.AN(\add_x_19_1/n184 ));
   XOR2X1TS U1368 (.Y(\addr_calc/fft_write_addr[2] ), 
	.B(n1454), 
	.A(FE_OCP_RBN1955_add_x_19_1_n187));
   OA21XLTS U1369 (.Y(\addr_calc/fft_read_addr[0] ), 
	.B0(\add_x_19_0/n191 ), 
	.A1(FE_OFN461_offset_0_), 
	.A0(FE_OFN517_addr_calc_fft_read_calc_count_0_));
   NOR3BX1TS U1370 (.Y(\data_cntl/N264 ), 
	.C(FE_OFN318_data_cntl_N95), 
	.B(FE_OFN330_data_to_fir), 
	.AN(n936));
   XOR2X1TS U1371 (.Y(\DP_OP_159_297_3515/n87 ), 
	.B(\add_x_22_4/n15 ), 
	.A(n1661));
   XOR2X4TS U1372 (.Y(n2593), 
	.B(n2366), 
	.A(\DP_OP_158_296_6262/n1998 ));
   XOR2XLTS U1373 (.Y(\DP_OP_159_297_3515/n556 ), 
	.B(n1964), 
	.A(\DP_OP_159_297_3515/n792 ));
   XNOR2X4TS U1374 (.Y(\addr_calc/fir_read_addr[21] ), 
	.B(n1569), 
	.A(n1568));
   NOR2XLTS U1375 (.Y(\DP_OP_158_296_6262/n1883 ), 
	.B(FE_OFN475_filesize_22_), 
	.A(\DP_OP_158_296_6262/n1891 ));
   NAND2X1TS U1376 (.Y(\DP_OP_159_297_3515/n646 ), 
	.B(\DP_OP_159_297_3515/n672 ), 
	.A(\DP_OP_159_297_3515/n648 ));
   XNOR2X1TS U1377 (.Y(\DP_OP_159_297_3515/n674 ), 
	.B(n2570), 
	.A(n2617));
   NOR2X4TS U1378 (.Y(\DP_OP_159_297_3515/n85 ), 
	.B(\DP_OP_159_297_3515/n87 ), 
	.A(\DP_OP_159_297_3515/n102 ));
   XOR2X4TS U1379 (.Y(\DP_OP_159_297_3515/n116 ), 
	.B(n2033), 
	.A(n1738));
   NAND2X2TS U1380 (.Y(\add_x_19_4/n185 ), 
	.B(FE_OCPUNCON1076_FE_OFN451_offset_2_), 
	.A(\addr_calc/iir_read_calc/count[2] ));
   AO22X1TS U1381 (.Y(n964), 
	.B1(\addr_calc/iir_read_calc/count[7] ), 
	.B0(FE_OFN93_n1192), 
	.A1(\addr_calc/iir_read_calc/counter/N50 ), 
	.A0(FE_OFN84_n2787));
   NOR2X1TS U1384 (.Y(\DP_OP_158_296_6262/n264 ), 
	.B(\DP_OP_158_296_6262/n266 ), 
	.A(\DP_OP_158_296_6262/n277 ));
   XOR2X1TS U1385 (.Y(\DP_OP_158_296_6262/n998 ), 
	.B(n1946), 
	.A(n1655));
   NAND2XLTS U1386 (.Y(n1734), 
	.B(\DP_OP_159_297_3515/n873 ), 
	.A(\DP_OP_159_297_3515/n1024 ));
   NAND2X1TS U1387 (.Y(\DP_OP_159_297_3515/n1024 ), 
	.B(\DP_OP_159_297_3515/n1025 ), 
	.A(n1788));
   CLKINVX2TS U1388 (.Y(n1787), 
	.A(FE_OFN519_DP_OP_159_297_3515_n1039));
   INVXLTS U1389 (.Y(n1455), 
	.A(\DP_OP_158_296_6262/n1959 ));
   XNOR2X4TS U1390 (.Y(\addr_calc/fir_read_addr[15] ), 
	.B(\add_x_19_2/n17 ), 
	.A(\add_x_19_2/n122 ));
   CLKXOR2X2TS U1391 (.Y(n2610), 
	.B(\DP_OP_159_297_3515/n878 ), 
	.A(\DP_OP_159_297_3515/n1057 ));
   NOR2X2TS U1392 (.Y(\DP_OP_159_297_3515/n1057 ), 
	.B(\DP_OP_159_297_3515/n879 ), 
	.A(\DP_OP_159_297_3515/n1063 ));
   OAI21X2TS U1393 (.Y(n1596), 
	.B0(\add_x_19_2/n82 ), 
	.A1(\add_x_19_2/n81 ), 
	.A0(\add_x_19_2/n83 ));
   CLKINVX6TS U1394 (.Y(n1788), 
	.A(FE_OFN519_DP_OP_159_297_3515_n1039));
   NAND2X4TS U1396 (.Y(\DP_OP_159_297_3515/n18 ), 
	.B(n1623), 
	.A(n1624));
   XNOR2X1TS U1397 (.Y(\DP_OP_158_296_6262/n1171 ), 
	.B(n2046), 
	.A(n1756));
   NAND2X6TS U1398 (.Y(\DP_OP_159_297_3515/n1026 ), 
	.B(FE_OFN491_filesize_9_), 
	.A(FE_OFN490_filesize_10_));
   AOI21X4TS U1399 (.Y(\add_x_19_1/n38 ), 
	.B0(n1546), 
	.A1(n2632), 
	.A0(\add_x_19_1/n43 ));
   NOR2X6TS U1401 (.Y(n1591), 
	.B(FE_OFN489_filesize_11_), 
	.A(FE_OFN490_filesize_10_));
   AO22X1TS U1403 (.Y(n981), 
	.B1(\addr_calc/iir_write_calc/count[21] ), 
	.B0(FE_OCPUNCON1572_n2812), 
	.A1(\addr_calc/iir_write_calc/counter/N64 ), 
	.A0(FE_OCPUNCON1883_n2813));
   XNOR2X1TS U1404 (.Y(\DP_OP_159_297_3515/n723 ), 
	.B(n2562), 
	.A(n2608));
   XOR2X1TS U1405 (.Y(n2608), 
	.B(\DP_OP_159_297_3515/n875 ), 
	.A(n1787));
   NAND2X1TS U1406 (.Y(\DP_OP_159_297_3515/n998 ), 
	.B(FE_OFN487_filesize_13_), 
	.A(FE_OFN486_filesize_14_));
   XOR2X1TS U1408 (.Y(n1653), 
	.B(n1838), 
	.A(\DP_OP_158_296_6262/n829 ));
   NOR2X1TS U1409 (.Y(\DP_OP_158_296_6262/n1950 ), 
	.B(\DP_OP_158_296_6262/n1951 ), 
	.A(n1693));
   INVX2TS U1410 (.Y(\DP_OP_158_296_6262/n1952 ), 
	.A(FE_OFN488_filesize_12_));
   INVX2TS U1411 (.Y(\DP_OP_158_296_6262/n1966 ), 
	.A(FE_OFN490_filesize_10_));
   NOR2X2TS U1413 (.Y(\DP_OP_158_296_6262/n1862 ), 
	.B(FE_OFN471_filesize_24_), 
	.A(FE_OFN470_filesize_25_));
   NOR2X4TS U1414 (.Y(\DP_OP_158_296_6262/n1840 ), 
	.B(\DP_OP_158_296_6262/n1841 ), 
	.A(FE_OCPUNCON1082_n2589));
   XNOR2X1TS U1415 (.Y(\DP_OP_158_296_6262/n933 ), 
	.B(FE_OFN275_addr_calc_fft_read_calc_count_29_), 
	.A(n1463));
   CLKINVX4TS U1417 (.Y(n1641), 
	.A(FE_OFN499_filesize_2_));
   INVX4TS U1420 (.Y(\DP_OP_158_296_6262/n841 ), 
	.A(\DP_OP_158_296_6262/n2048 ));
   XNOR2X1TS U1421 (.Y(n1459), 
	.B(\add_x_22_0/n49 ), 
	.A(\DP_OP_158_296_6262/n2048 ));
   NOR2X1TS U1424 (.Y(\DP_OP_158_296_6262/n1077 ), 
	.B(\DP_OP_158_296_6262/n1079 ), 
	.A(n1459));
   AO22X1TS U1425 (.Y(n1121), 
	.B1(n1872), 
	.B0(FE_OCPUNCON1083_n2805), 
	.A1(\addr_calc/fir_write_calc/counter/N52 ), 
	.A0(FE_OFN547_n2803));
   OAI2BB1X1TS U1427 (.Y(n1110), 
	.B0(n1618), 
	.A1N(FE_OCPUNCON1087_n2805), 
	.A0N(\addr_calc/fir_write_calc/count[20] ));
   XOR2X4TS U1428 (.Y(n2625), 
	.B(n2341), 
	.A(\DP_OP_159_297_3515/n892 ));
   CLKINVX4TS U1429 (.Y(n783), 
	.A(\addr_calc/fft_read_calc/counter/N38 ));
   XOR2X4TS U1430 (.Y(\DP_OP_158_296_6262/n962 ), 
	.B(n1943), 
	.A(FE_OCPN1947_n1149));
   NOR2X4TS U1431 (.Y(n2807), 
	.B(n1461), 
	.A(n1696));
   XNOR2X1TS U1432 (.Y(\DP_OP_158_296_6262/n68 ), 
	.B(FE_OFN243_addr_calc_fir_read_calc_count_27_), 
	.A(n1149));
   AND2X8TS U1437 (.Y(n1461), 
	.B(n1715), 
	.A(n1716));
   NOR2X2TS U1438 (.Y(\DP_OP_158_296_6262/n1881 ), 
	.B(\DP_OP_158_296_6262/n1882 ), 
	.A(n1717));
   XOR2X2TS U1439 (.Y(\DP_OP_159_297_3515/n131 ), 
	.B(\add_x_22_4/n30 ), 
	.A(\DP_OP_159_297_3515/n792 ));
   AO22X1TS U1440 (.Y(n1088), 
	.B1(FE_OFN63_n2809), 
	.B0(\addr_calc/fir_read_calc/count[10] ), 
	.A1(\addr_calc/fir_read_calc/counter/N53 ), 
	.A0(FE_OFN54_n2807));
   AO22X1TS U1441 (.Y(n1077), 
	.B1(FE_OFN66_n2809), 
	.B0(\addr_calc/fir_read_calc/count[21] ), 
	.A1(\addr_calc/fir_read_calc/counter/N64 ), 
	.A0(FE_OFN56_n2807));
   NOR2X1TS U1442 (.Y(\DP_OP_158_296_6262/n1109 ), 
	.B(\DP_OP_158_296_6262/n1124 ), 
	.A(\DP_OP_158_296_6262/n1111 ));
   XNOR2X1TS U1443 (.Y(\DP_OP_158_296_6262/n1111 ), 
	.B(FE_OFN287_addr_calc_fft_read_calc_count_17_), 
	.A(n1729));
   NAND2X1TS U1444 (.Y(\add_x_22_1/n3 ), 
	.B(\add_x_22_1/n59 ), 
	.A(\add_x_22_1/n4 ));
   XNOR2X1TS U1445 (.Y(\DP_OP_158_296_6262/n54 ), 
	.B(n1775), 
	.A(n1871));
   OAI21X4TS U1446 (.Y(\add_x_19_2/n134 ), 
	.B0(\add_x_19_2/n136 ), 
	.A1(\add_x_19_2/n135 ), 
	.A0(\add_x_19_2/n156 ));
   NOR2X1TS U1447 (.Y(\DP_OP_158_296_6262/n1964 ), 
	.B(\DP_OP_158_296_6262/n1965 ), 
	.A(n1693));
   AND2X2TS U1448 (.Y(n1462), 
	.B(\DP_OP_158_296_6262/n1869 ), 
	.A(\DP_OP_158_296_6262/n1791 ));
   INVX6TS U1449 (.Y(n1717), 
	.A(n1677));
   AO22X1TS U1450 (.Y(n954), 
	.B1(\addr_calc/iir_read_calc/count[17] ), 
	.B0(FE_OFN90_n1192), 
	.A1(\addr_calc/iir_read_calc/counter/N60 ), 
	.A0(FE_OFN78_n2787));
   XNOR2X2TS U1451 (.Y(\addr_calc/fft_write_addr[15] ), 
	.B(\add_x_19_1/n17 ), 
	.A(\add_x_19_1/n122 ));
   XNOR2X1TS U1452 (.Y(\DP_OP_158_296_6262/n148 ), 
	.B(\addr_calc/fir_read_calc/count[22] ), 
	.A(n1652));
   AO22X1TS U1453 (.Y(n1049), 
	.B1(n1924), 
	.B0(FE_OFN20_n2797), 
	.A1(\addr_calc/fft_write_calc/counter/N60 ), 
	.A0(FE_OFN29_n2795));
   AO22X1TS U1454 (.Y(n1050), 
	.B1(n2567), 
	.B0(FE_OFN19_n2797), 
	.A1(\addr_calc/fft_write_calc/counter/N59 ), 
	.A0(FE_OFN28_n2795));
   XOR2X1TS U1455 (.Y(n1471), 
	.B(FE_OFN278_addr_calc_fft_read_calc_count_30_), 
	.A(\DP_OP_158_296_6262/n829 ));
   NOR2X2TS U1456 (.Y(\DP_OP_158_296_6262/n1847 ), 
	.B(\DP_OP_158_296_6262/n1848 ), 
	.A(FE_OCPUNCON1082_n2589));
   XOR2X4TS U1457 (.Y(n1463), 
	.B(n1464), 
	.A(\DP_OP_158_296_6262/n1840 ));
   NOR2X4TS U1458 (.Y(\DP_OP_158_296_6262/n1791 ), 
	.B(\DP_OP_158_296_6262/n1877 ), 
	.A(\DP_OP_158_296_6262/n1903 ));
   NAND2X2TS U1459 (.Y(\DP_OP_158_296_6262/n1877 ), 
	.B(\DP_OP_158_296_6262/n1878 ), 
	.A(\DP_OP_158_296_6262/n1890 ));
   NAND2X1TS U1460 (.Y(\DP_OP_158_296_6262/n1848 ), 
	.B(\DP_OP_158_296_6262/n1849 ), 
	.A(FE_OFN113_DP_OP_158_296_6262_n1791));
   AO22X4TS U1461 (.Y(n1061), 
	.B1(n1479), 
	.B0(FE_OFN26_n2797), 
	.A1(\addr_calc/fft_write_calc/counter/N48 ), 
	.A0(FE_OFN35_n2795));
   XNOR2X4TS U1463 (.Y(\addr_calc/fft_write_addr[23] ), 
	.B(\add_x_19_1/n9 ), 
	.A(\add_x_19_1/n80 ));
   OR2X4TS U1464 (.Y(n1693), 
	.B(\DP_OP_158_296_6262/n1987 ), 
	.A(\DP_OP_158_296_6262/n2011 ));
   CLKINVX2TS U1465 (.Y(\DP_OP_159_297_3515/n876 ), 
	.A(FE_OFN492_filesize_8_));
   XNOR2X1TS U1466 (.Y(\DP_OP_159_297_3515/n650 ), 
	.B(n1951), 
	.A(n2615));
   NOR2X4TS U1467 (.Y(\add_x_19_2/n162 ), 
	.B(\addr_calc/fir_read_calc/count[7] ), 
	.A(FE_OCP_RBN1841_offset_7_));
   NAND2X2TS U1468 (.Y(\add_x_19_2/n163 ), 
	.B(FE_OCP_RBN1841_offset_7_), 
	.A(\addr_calc/fir_read_calc/count[7] ));
   NAND2X2TS U1471 (.Y(\DP_OP_158_296_6262/n958 ), 
	.B(\DP_OP_158_296_6262/n996 ), 
	.A(\DP_OP_158_296_6262/n960 ));
   NOR2X1TS U1472 (.Y(\DP_OP_158_296_6262/n1895 ), 
	.B(FE_OCPUNCON1081_n2589), 
	.A(\DP_OP_158_296_6262/n1896 ));
   NOR2X4TS U1473 (.Y(\DP_OP_158_296_6262/n62 ), 
	.B(\DP_OP_158_296_6262/n64 ), 
	.A(\DP_OP_158_296_6262/n129 ));
   NOR2X6TS U1474 (.Y(n1736), 
	.B(\DP_OP_158_296_6262/n1854 ), 
	.A(FE_OCPUNCON1567_n1717));
   AOI21X4TS U1476 (.Y(\add_x_19_2/n60 ), 
	.B0(\add_x_19_2/n62 ), 
	.A1(\add_x_19_2/n61 ), 
	.A0(\add_x_19_2/n69 ));
   OAI21X2TS U1477 (.Y(\add_x_19_2/n92 ), 
	.B0(\add_x_19_2/n94 ), 
	.A1(\add_x_19_2/n93 ), 
	.A0(FE_OFN526_add_x_19_2_n113));
   NOR2X4TS U1478 (.Y(\DP_OP_158_296_6262/n956 ), 
	.B(\DP_OP_158_296_6262/n958 ), 
	.A(\DP_OP_158_296_6262/n1023 ));
   NAND2X2TS U1479 (.Y(\DP_OP_158_296_6262/n1023 ), 
	.B(\DP_OP_158_296_6262/n1053 ), 
	.A(\DP_OP_158_296_6262/n1025 ));
   NOR2X1TS U1481 (.Y(\DP_OP_158_296_6262/n1860 ), 
	.B(\DP_OP_158_296_6262/n1861 ), 
	.A(FE_OCPUNCON1082_n2589));
   OAI2BB2XLTS U1483 (.Y(n989), 
	.B1(\add_x_22_5/n71 ), 
	.B0(n1740), 
	.A1N(\addr_calc/iir_write_calc/counter/N56 ), 
	.A0N(FE_OCPUNCON1879_n2813));
   XNOR2X1TS U1484 (.Y(\DP_OP_159_297_3515/n714 ), 
	.B(n1940), 
	.A(n2621));
   XOR2X4TS U1487 (.Y(n2594), 
	.B(FE_OFN482_filesize_16_), 
	.A(n1717));
   XNOR2X4TS U1489 (.Y(\addr_calc/fft_write_addr[27] ), 
	.B(\add_x_19_1/n5 ), 
	.A(\add_x_19_1/n57 ));
   NOR2X2TS U1490 (.Y(\DP_OP_158_296_6262/n1890 ), 
	.B(FE_OFN476_filesize_21_), 
	.A(FE_OFN477_filesize_20_));
   NOR2X1TS U1493 (.Y(n1642), 
	.B(\DP_OP_158_296_6262/n1903 ), 
	.A(FE_OCPUNCON1081_n2589));
   NOR2X4TS U1495 (.Y(\DP_OP_158_296_6262/n1973 ), 
	.B(FE_OFN491_filesize_9_), 
	.A(FE_OFN492_filesize_8_));
   INVXLTS U1496 (.Y(\DP_OP_158_296_6262/n1946 ), 
	.A(\DP_OP_158_296_6262/n1945 ));
   CLKINVX3TS U1498 (.Y(n2006), 
	.A(n2005));
   INVX2TS U1499 (.Y(\DP_OP_158_296_6262/n1911 ), 
	.A(FE_OFN479_filesize_18_));
   CLKINVX2TS U1501 (.Y(n1918), 
	.A(n1917));
   INVX2TS U1502 (.Y(n1989), 
	.A(\addr_calc/fir_write_calc/count[2] ));
   INVX2TS U1503 (.Y(n2057), 
	.A(FE_OFN517_addr_calc_fft_read_calc_count_0_));
   INVX2TS U1504 (.Y(n2330), 
	.A(FE_OFN466_filesize_28_));
   INVX2TS U1505 (.Y(n1533), 
	.A(\add_x_19_5/n36 ));
   AND2X2TS U1506 (.Y(n1465), 
	.B(\add_x_19_0/n56 ), 
	.A(\add_x_19_0/n196 ));
   AND2X2TS U1507 (.Y(n1466), 
	.B(\add_x_19_4/n79 ), 
	.A(\add_x_19_4/n200 ));
   INVXLTS U1508 (.Y(\DP_OP_159_297_3515/n869 ), 
	.A(FE_OFN483_filesize_15_));
   CLKAND2X2TS U1509 (.Y(n1467), 
	.B(\add_x_19_4/n67 ), 
	.A(\add_x_19_4/n199 ));
   OR3X1TS U1510 (.Y(n1468), 
	.C(n1861), 
	.B(n2790), 
	.A(FE_OFN314_data_cntl_N159));
   INVX2TS U1512 (.Y(\DP_OP_158_296_6262/n1869 ), 
	.A(FE_OFN471_filesize_24_));
   INVXLTS U1513 (.Y(n2367), 
	.A(\DP_OP_158_296_6262/n1966 ));
   INVXLTS U1514 (.Y(\DP_OP_159_297_3515/n870 ), 
	.A(FE_OFN485_filesize_14_));
   INVXLTS U1515 (.Y(n2368), 
	.A(\DP_OP_158_296_6262/n1952 ));
   CLKINVX12TS U1517 (.Y(n1677), 
	.A(FE_OCPUNCON1082_n2589));
   XNOR2X4TS U1518 (.Y(n1469), 
	.B(n2365), 
	.A(\DP_OP_158_296_6262/n1978 ));
   INVX2TS U1519 (.Y(\add_x_19_3/n123 ), 
	.A(n1545));
   CLKAND2X2TS U1520 (.Y(n1470), 
	.B(\add_x_19_3/n46 ), 
	.A(\add_x_19_3/n72 ));
   INVX2TS U1521 (.Y(n2371), 
	.A(\DP_OP_159_297_3515/n880 ));
   INVX2TS U1524 (.Y(n1901), 
	.A(\addr_calc/iir_read_calc/count[3] ));
   INVX2TS U1525 (.Y(n1925), 
	.A(\addr_calc/iir_read_calc/count[25] ));
   INVX2TS U1527 (.Y(n1897), 
	.A(\addr_calc/fir_read_calc/count[10] ));
   INVX2TS U1528 (.Y(\addr_calc/fir_write_calc/counter/N43 ), 
	.A(\addr_calc/fir_write_calc/count[0] ));
   NAND2X1TS U1561 (.Y(\DP_OP_159_297_3515/n1052 ), 
	.B(FE_OFN495_filesize_5_), 
	.A(FE_OFN494_filesize_6_));
   INVXLTS U1562 (.Y(\DP_OP_159_297_3515/n878 ), 
	.A(FE_OFN494_filesize_6_));
   INVXLTS U1563 (.Y(\DP_OP_159_297_3515/n950 ), 
	.A(FE_OFN476_filesize_21_));
   NAND2X1TS U1564 (.Y(\DP_OP_159_297_3515/n943 ), 
	.B(FE_OFN474_filesize_22_), 
	.A(FE_OFN476_filesize_21_));
   OAI21XLTS U1568 (.Y(n1536), 
	.B0(\add_x_19_5/n124 ), 
	.A1(\add_x_19_5/n123 ), 
	.A0(\add_x_19_5/n125 ));
   CLKINVX1TS U1570 (.Y(\add_x_19_1/n200 ), 
	.A(\add_x_19_1/n78 ));
   AO21X4TS U1571 (.Y(\add_x_19_5/n35 ), 
	.B0(n1534), 
	.A1(FE_OFN531_add_x_19_5_n43), 
	.A0(n1532));
   XNOR2X4TS U1572 (.Y(\addr_calc/iir_write_addr[31] ), 
	.B(\add_x_19_5/n1 ), 
	.A(\add_x_19_5/n35 ));
   OAI21X2TS U1573 (.Y(\add_x_19_5/n73 ), 
	.B0(\add_x_19_5/n75 ), 
	.A1(\add_x_19_5/n74 ), 
	.A0(\add_x_19_5/n94 ));
   NAND2X2TS U1574 (.Y(\add_x_19_0/n132 ), 
	.B(FE_OFN413_offset_12_), 
	.A(n2046));
   AOI21X1TS U1575 (.Y(\add_x_19_5/n45 ), 
	.B0(\add_x_19_5/n47 ), 
	.A1(\add_x_19_5/n46 ), 
	.A0(\add_x_19_5/n73 ));
   NAND2X1TS U1576 (.Y(\add_x_19_5/n44 ), 
	.B(\add_x_19_5/n46 ), 
	.A(\add_x_19_5/n72 ));
   OAI21X1TS U1577 (.Y(\add_x_19_5/n43 ), 
	.B0(\add_x_19_5/n45 ), 
	.A1(\add_x_19_5/n44 ), 
	.A0(\add_x_19_5/n113 ));
   OAI21X4TS U1578 (.Y(\add_x_19_5/n134 ), 
	.B0(\add_x_19_5/n136 ), 
	.A1(\add_x_19_5/n135 ), 
	.A0(\add_x_19_5/n156 ));
   XNOR2X2TS U1580 (.Y(\addr_calc/iir_write_addr[15] ), 
	.B(n1537), 
	.A(n1536));
   INVX1TS U1581 (.Y(\add_x_22_2/n98 ), 
	.A(\addr_calc/fir_read_calc/count[7] ));
   CLKINVX1TS U1582 (.Y(\add_x_19_2/n216 ), 
	.A(\add_x_19_2/n162 ));
   INVX3TS U1583 (.Y(\add_x_19_2/n156 ), 
	.A(FE_OFN122_add_x_19_2_n157));
   OAI21X4TS U1584 (.Y(\add_x_19_0/n115 ), 
	.B0(\add_x_19_0/n117 ), 
	.A1(n1539), 
	.A0(\add_x_19_0/n136 ));
   NOR2X8TS U1585 (.Y(\add_x_19_0/n114 ), 
	.B(n1539), 
	.A(\add_x_19_0/n135 ));
   NAND2X2TS U1586 (.Y(n1539), 
	.B(\add_x_19_0/n126 ), 
	.A(\add_x_19_0/n118 ));
   NAND2X6TS U1587 (.Y(\add_x_19_3/n191 ), 
	.B(FE_OFN252_addr_calc_fir_write_calc_count_0_), 
	.A(FE_OFN461_offset_0_));
   NAND2X4TS U1588 (.Y(\add_x_19_3/n185 ), 
	.B(FE_OFN452_offset_2_), 
	.A(n1990));
   NOR2X2TS U1589 (.Y(\add_x_19_2/n144 ), 
	.B(FE_OCPUNCON653_FE_OFN418_offset_10_), 
	.A(n1540));
   NAND2X2TS U1590 (.Y(\add_x_19_2/n145 ), 
	.B(FE_OCPUNCON653_FE_OFN418_offset_10_), 
	.A(n1540));
   XNOR2X1TS U1591 (.Y(\DP_OP_158_296_6262/n297 ), 
	.B(n1540), 
	.A(n1656));
   INVX1TS U1592 (.Y(\add_x_19_2/n143 ), 
	.A(\add_x_19_2/n145 ));
   INVX6TS U1593 (.Y(\add_x_19_2/n112 ), 
	.A(FE_OFN526_add_x_19_2_n113));
   XNOR2X1TS U1595 (.Y(n1543), 
	.B(\addr_calc/fft_read_calc/count[31] ), 
	.A(\add_x_22_0/n1 ));
   OAI2BB1X1TS U1596 (.Y(n1035), 
	.B0(n1542), 
	.A1N(FE_OFN15_n2794), 
	.A0N(\addr_calc/fft_read_calc/count[31] ));
   OAI21X4TS U1598 (.Y(\add_x_19_3/n169 ), 
	.B0(\add_x_19_3/n171 ), 
	.A1(\add_x_19_3/n170 ), 
	.A0(\add_x_19_3/n176 ));
   OAI21X4TS U1600 (.Y(\add_x_19_3/n187 ), 
	.B0(\add_x_19_3/n189 ), 
	.A1(\add_x_19_3/n191 ), 
	.A0(\add_x_19_3/n188 ));
   OAI21X2TS U1601 (.Y(\add_x_19_2/n150 ), 
	.B0(\add_x_19_2/n152 ), 
	.A1(\add_x_19_2/n155 ), 
	.A0(\add_x_19_2/n151 ));
   AOI21X2TS U1602 (.Y(\add_x_19_2/n45 ), 
	.B0(\add_x_19_2/n47 ), 
	.A1(\add_x_19_2/n46 ), 
	.A0(\add_x_19_2/n73 ));
   NAND2X4TS U1603 (.Y(\add_x_19_5/n116 ), 
	.B(\add_x_19_5/n126 ), 
	.A(\add_x_19_5/n118 ));
   NOR2X1TS U1604 (.Y(n1547), 
	.B(\add_x_19_2/n184 ), 
	.A(\add_x_19_2/n181 ));
   AOI21X4TS U1607 (.Y(\add_x_19_5/n113 ), 
	.B0(FE_OFN140_add_x_19_5_n115), 
	.A1(FE_OFN522_add_x_19_5_n114), 
	.A0(FE_OFN129_add_x_19_5_n157));
   OAI21X2TS U1608 (.Y(\add_x_19_5/n92 ), 
	.B0(\add_x_19_5/n94 ), 
	.A1(\add_x_19_5/n93 ), 
	.A0(\add_x_19_5/n113 ));
   NOR2X6TS U1609 (.Y(\add_x_19_3/n120 ), 
	.B(FE_OFN400_offset_15_), 
	.A(n1883));
   NOR2X4TS U1610 (.Y(\add_x_19_3/n118 ), 
	.B(\add_x_19_3/n120 ), 
	.A(\add_x_19_3/n123 ));
   INVX1TS U1613 (.Y(\add_x_19_0/n196 ), 
	.A(\add_x_19_0/n55 ));
   NOR2X2TS U1614 (.Y(n1549), 
	.B(\add_x_19_4/n120 ), 
	.A(\add_x_19_4/n123 ));
   NAND2X2TS U1615 (.Y(n1567), 
	.B(n1549), 
	.A(\add_x_19_4/n126 ));
   NOR2X8TS U1616 (.Y(\add_x_19_1/n170 ), 
	.B(\addr_calc/fft_write_calc/count[5] ), 
	.A(FE_OCP_RBN1493_offset_5_));
   NOR2X4TS U1617 (.Y(\add_x_19_3/n126 ), 
	.B(\add_x_19_3/n131 ), 
	.A(\add_x_19_3/n128 ));
   NOR2X6TS U1618 (.Y(\add_x_19_3/n184 ), 
	.B(FE_OFN452_offset_2_), 
	.A(n1990));
   NOR2X6TS U1620 (.Y(\add_x_19_0/n128 ), 
	.B(n1967), 
	.A(FE_OCPUNCON1943_FE_OFN407_offset_13_));
   NAND2X2TS U1621 (.Y(\add_x_19_3/n116 ), 
	.B(\add_x_19_3/n126 ), 
	.A(\add_x_19_3/n118 ));
   AOI2BB1X4TS U1622 (.Y(\addr_calc/fft_write_addr[31] ), 
	.B0(n1551), 
	.A1N(n1550), 
	.A0N(\add_x_19_1/n38 ));
   INVX2TS U1625 (.Y(\add_x_19_1/n71 ), 
	.A(\add_x_19_1/n73 ));
   INVX2TS U1626 (.Y(\add_x_19_1/n70 ), 
	.A(\add_x_19_1/n72 ));
   AOI21X4TS U1627 (.Y(\add_x_19_5/n102 ), 
	.B0(\add_x_19_5/n104 ), 
	.A1(\add_x_19_5/n103 ), 
	.A0(\add_x_19_5/n112 ));
   INVX1TS U1628 (.Y(\add_x_19_1/n196 ), 
	.A(\add_x_19_1/n55 ));
   INVX1TS U1629 (.Y(\add_x_19_5/n204 ), 
	.A(\add_x_19_5/n97 ));
   AOI21X4TS U1632 (.Y(\add_x_19_0/n113 ), 
	.B0(\add_x_19_0/n115 ), 
	.A1(\add_x_19_0/n114 ), 
	.A0(FE_OFN139_add_x_19_0_n157));
   INVX4TS U1633 (.Y(\add_x_19_0/n156 ), 
	.A(FE_OFN139_add_x_19_0_n157));
   OAI21X4TS U1634 (.Y(\add_x_19_0/n43 ), 
	.B0(\add_x_19_0/n45 ), 
	.A1(\add_x_19_0/n44 ), 
	.A0(FE_OFN528_add_x_19_0_n113));
   OAI21X4TS U1637 (.Y(\add_x_19_0/n80 ), 
	.B0(\add_x_19_0/n82 ), 
	.A1(\add_x_19_0/n81 ), 
	.A0(\add_x_19_0/n83 ));
   XOR2X4TS U1638 (.Y(\addr_calc/fft_read_addr[23] ), 
	.B(n1561), 
	.A(\add_x_19_0/n80 ));
   OR2X1TS U1639 (.Y(n1560), 
	.B(FE_OFN337_offset_31_), 
	.A(FE_OFN261_addr_calc_fir_read_calc_count_31_));
   INVX1TS U1640 (.Y(\add_x_19_0/n200 ), 
	.A(\add_x_19_0/n78 ));
   AND2X6TS U1641 (.Y(n1561), 
	.B(\add_x_19_0/n79 ), 
	.A(\add_x_19_0/n200 ));
   NOR2X6TS U1642 (.Y(\add_x_19_3/n162 ), 
	.B(FE_OCPUNCON1278_offset_7_), 
	.A(\addr_calc/fir_write_calc/count[7] ));
   INVX1TS U1644 (.Y(\DP_OP_159_297_3515/n901 ), 
	.A(\DP_OP_159_297_3515/n902 ));
   NAND2X2TS U1645 (.Y(\DP_OP_159_297_3515/n899 ), 
	.B(\DP_OP_159_297_3515/n900 ), 
	.A(FE_OCPUNCON1566_n1789));
   XOR2X4TS U1646 (.Y(n2613), 
	.B(FE_OFN464_filesize_29_), 
	.A(\DP_OP_159_297_3515/n899 ));
   XNOR2X1TS U1647 (.Y(\DP_OP_159_297_3515/n541 ), 
	.B(n2051), 
	.A(n1738));
   XNOR2XLTS U1648 (.Y(\DP_OP_159_297_3515/n569 ), 
	.B(n2579), 
	.A(n1703));
   XOR2X1TS U1649 (.Y(\DP_OP_159_297_3515/n582 ), 
	.B(n1961), 
	.A(n1699));
   XOR2X2TS U1650 (.Y(\DP_OP_159_297_3515/n476 ), 
	.B(\addr_calc/iir_write_calc/count[28] ), 
	.A(\DP_OP_159_297_3515/n1138 ));
   XOR2X1TS U1651 (.Y(\DP_OP_159_297_3515/n527 ), 
	.B(n1968), 
	.A(n1732));
   XNOR2X1TS U1652 (.Y(\DP_OP_159_297_3515/n512 ), 
	.B(n2573), 
	.A(n1661));
   NOR2X1TS U1653 (.Y(\DP_OP_159_297_3515/n539 ), 
	.B(\DP_OP_159_297_3515/n541 ), 
	.A(\DP_OP_159_297_3515/n556 ));
   NOR2X1TS U1654 (.Y(\DP_OP_159_297_3515/n567 ), 
	.B(\DP_OP_159_297_3515/n569 ), 
	.A(\DP_OP_159_297_3515/n582 ));
   NOR2X1TS U1655 (.Y(\DP_OP_159_297_3515/n474 ), 
	.B(\DP_OP_159_297_3515/n495 ), 
	.A(\DP_OP_159_297_3515/n476 ));
   NOR2X1TS U1656 (.Y(\DP_OP_159_297_3515/n510 ), 
	.B(\DP_OP_159_297_3515/n527 ), 
	.A(\DP_OP_159_297_3515/n512 ));
   NAND2X2TS U1657 (.Y(\DP_OP_159_297_3515/n443 ), 
	.B(n1563), 
	.A(n1564));
   NAND2X1TS U1658 (.Y(\DP_OP_159_297_3515/n537 ), 
	.B(\DP_OP_159_297_3515/n539 ), 
	.A(\DP_OP_159_297_3515/n567 ));
   NAND2X2TS U1659 (.Y(\DP_OP_159_297_3515/n472 ), 
	.B(\DP_OP_159_297_3515/n474 ), 
	.A(\DP_OP_159_297_3515/n510 ));
   NOR2X2TS U1660 (.Y(\DP_OP_159_297_3515/n428 ), 
	.B(\DP_OP_159_297_3515/n430 ), 
	.A(\DP_OP_159_297_3515/n443 ));
   NOR2X2TS U1661 (.Y(\DP_OP_159_297_3515/n470 ), 
	.B(\DP_OP_159_297_3515/n537 ), 
	.A(\DP_OP_159_297_3515/n472 ));
   AND2X6TS U1662 (.Y(n1779), 
	.B(\DP_OP_159_297_3515/n428 ), 
	.A(\DP_OP_159_297_3515/n470 ));
   OAI2BB1X1TS U1664 (.Y(n986), 
	.B0(n1565), 
	.A1N(FE_OCPUNCON1570_n2812), 
	.A0N(n1951));
   OAI21X4TS U1668 (.Y(\add_x_19_4/n92 ), 
	.B0(\add_x_19_4/n94 ), 
	.A1(\add_x_19_4/n93 ), 
	.A0(FE_OFN527_add_x_19_4_n113));
   INVX6TS U1671 (.Y(\add_x_19_4/n112 ), 
	.A(FE_OFN527_add_x_19_4_n113));
   OAI21X2TS U1673 (.Y(\add_x_19_4/n80 ), 
	.B0(\add_x_19_4/n82 ), 
	.A1(\add_x_19_4/n81 ), 
	.A0(\add_x_19_4/n83 ));
   OAI21X4TS U1674 (.Y(\add_x_19_3/n150 ), 
	.B0(\add_x_19_3/n152 ), 
	.A1(\add_x_19_3/n151 ), 
	.A0(\add_x_19_3/n155 ));
   CLKINVX1TS U1675 (.Y(\add_x_19_4/n200 ), 
	.A(\add_x_19_4/n78 ));
   XOR2X4TS U1676 (.Y(\addr_calc/iir_read_addr[23] ), 
	.B(n1466), 
	.A(\add_x_19_4/n80 ));
   NAND2BX1TS U1678 (.Y(n1570), 
	.B(FE_OFN81_n2787), 
	.AN(n1571));
   OAI2BB1X1TS U1679 (.Y(n945), 
	.B0(n1570), 
	.A1N(FE_OFN88_n2654), 
	.A0N(n1572));
   INVX1TS U1680 (.Y(\add_x_19_5/n200 ), 
	.A(\add_x_19_5/n78 ));
   OAI21X4TS U1682 (.Y(\add_x_19_3/n127 ), 
	.B0(\add_x_19_3/n129 ), 
	.A1(\add_x_19_3/n128 ), 
	.A0(\add_x_19_3/n132 ));
   NAND2BX1TS U1683 (.Y(n1573), 
	.B(FE_OCPUNCON1881_n2813), 
	.AN(n1574));
   OAI2BB1X1TS U1684 (.Y(n987), 
	.B0(n1573), 
	.A1N(FE_OCPUNCON1568_n2812), 
	.A0N(\addr_calc/iir_write_calc/count[15] ));
   NAND2BX1TS U1685 (.Y(n1576), 
	.B(FE_OFN81_n2787), 
	.AN(n1577));
   OAI2BB1X1TS U1686 (.Y(n944), 
	.B0(n1576), 
	.A1N(FE_OFN88_n2654), 
	.A0N(\addr_calc/iir_read_calc/count[27] ));
   OR2X2TS U1691 (.Y(n1586), 
	.B(FE_OFN340_offset_31_), 
	.A(FE_OFN234_addr_calc_iir_read_calc_count_31_));
   NOR2X2TS U1692 (.Y(n1587), 
	.B(\add_x_19_0/n184 ), 
	.A(\add_x_19_0/n181 ));
   AOI21X4TS U1693 (.Y(\add_x_19_0/n178 ), 
	.B0(n1588), 
	.A1(n1587), 
	.A0(\add_x_19_0/n187 ));
   OR2X2TS U1694 (.Y(n1590), 
	.B(FE_OFN340_offset_31_), 
	.A(FE_OFN240_addr_calc_iir_write_calc_count_31_));
   NOR2X4TS U1695 (.Y(n1592), 
	.B(\add_x_19_3/n116 ), 
	.A(\add_x_19_3/n135 ));
   AOI21X4TS U1696 (.Y(\add_x_19_3/n113 ), 
	.B0(n1593), 
	.A1(FE_OFN521_n1592), 
	.A0(FE_OFN525_add_x_19_3_n157));
   OAI21X4TS U1697 (.Y(n1593), 
	.B0(n1594), 
	.A1(\add_x_19_3/n116 ), 
	.A0(\add_x_19_3/n136 ));
   CLKINVX1TS U1699 (.Y(\add_x_19_3/n200 ), 
	.A(\add_x_19_3/n78 ));
   OAI21X2TS U1700 (.Y(\add_x_19_3/n80 ), 
	.B0(\add_x_19_3/n82 ), 
	.A1(\add_x_19_3/n81 ), 
	.A0(\add_x_19_3/n83 ));
   AOI21X2TS U1701 (.Y(\add_x_19_2/n83 ), 
	.B0(\add_x_19_2/n85 ), 
	.A1(\add_x_19_2/n84 ), 
	.A0(\add_x_19_2/n92 ));
   NOR2X1TS U1702 (.Y(\DP_OP_158_296_6262/n1850 ), 
	.B(FE_OFN468_filesize_26_), 
	.A(FE_OFN467_filesize_27_));
   NAND2X2TS U1703 (.Y(\DP_OP_158_296_6262/n1792 ), 
	.B(\DP_OP_158_296_6262/n1850 ), 
	.A(\DP_OP_158_296_6262/n1862 ));
   XOR2X1TS U1704 (.Y(n1598), 
	.B(\addr_calc/fft_read_calc/count[2] ), 
	.A(n2596));
   XOR2X1TS U1705 (.Y(n1601), 
	.B(FE_OFN264_addr_calc_fft_read_calc_count_4_), 
	.A(\DP_OP_158_296_6262/n855 ));
   XOR2X1TS U1706 (.Y(n1600), 
	.B(n1978), 
	.A(FE_OFN75_n2599));
   XOR2X1TS U1707 (.Y(n1599), 
	.B(FE_OFN225_addr_calc_fft_read_calc_count_6_), 
	.A(n2593));
   XNOR2X1TS U1708 (.Y(\DP_OP_158_296_6262/n1180 ), 
	.B(n1970), 
	.A(n1660));
   XOR2X1TS U1709 (.Y(\DP_OP_158_296_6262/n1079 ), 
	.B(n1955), 
	.A(n1654));
   XNOR2X1TS U1710 (.Y(\DP_OP_158_296_6262/n948 ), 
	.B(\addr_calc/fft_read_calc/count[28] ), 
	.A(n1775));
   XOR2X4TS U1711 (.Y(\DP_OP_158_296_6262/n1013 ), 
	.B(n2037), 
	.A(FE_OCPN1732_n1718));
   XOR2X1TS U1712 (.Y(\DP_OP_158_296_6262/n981 ), 
	.B(\add_x_22_0/n15 ), 
	.A(\DP_OP_158_296_6262/n833 ));
   XNOR2X1TS U1713 (.Y(\DP_OP_158_296_6262/n1068 ), 
	.B(n2572), 
	.A(n1776));
   NOR2X1TS U1714 (.Y(\DP_OP_158_296_6262/n1241 ), 
	.B(\DP_OP_158_296_6262/n1259 ), 
	.A(\DP_OP_158_296_6262/n1243 ));
   NOR2X1TS U1715 (.Y(\DP_OP_158_296_6262/n1214 ), 
	.B(\DP_OP_158_296_6262/n1223 ), 
	.A(\DP_OP_158_296_6262/n1216 ));
   NOR2X1TS U1716 (.Y(\DP_OP_158_296_6262/n1198 ), 
	.B(\DP_OP_158_296_6262/n1209 ), 
	.A(\DP_OP_158_296_6262/n1200 ));
   NOR2X1TS U1717 (.Y(\DP_OP_158_296_6262/n1178 ), 
	.B(\DP_OP_158_296_6262/n1180 ), 
	.A(\DP_OP_158_296_6262/n1191 ));
   NOR2X1TS U1718 (.Y(\DP_OP_158_296_6262/n1134 ), 
	.B(\DP_OP_158_296_6262/n1136 ), 
	.A(\DP_OP_158_296_6262/n1149 ));
   NOR2X1TS U1719 (.Y(\DP_OP_158_296_6262/n931 ), 
	.B(\DP_OP_158_296_6262/n948 ), 
	.A(\DP_OP_158_296_6262/n933 ));
   NOR2X2TS U1720 (.Y(\DP_OP_158_296_6262/n960 ), 
	.B(\DP_OP_158_296_6262/n962 ), 
	.A(\DP_OP_158_296_6262/n981 ));
   NOR2X1TS U1721 (.Y(\DP_OP_158_296_6262/n1025 ), 
	.B(\DP_OP_158_296_6262/n1027 ), 
	.A(\DP_OP_158_296_6262/n1042 ));
   NOR2X1TS U1722 (.Y(\DP_OP_158_296_6262/n1053 ), 
	.B(\DP_OP_158_296_6262/n1055 ), 
	.A(\DP_OP_158_296_6262/n1068 ));
   NAND2X4TS U1723 (.Y(\DP_OP_158_296_6262/n1212 ), 
	.B(\DP_OP_158_296_6262/n1241 ), 
	.A(\DP_OP_158_296_6262/n1214 ));
   NAND2X1TS U1724 (.Y(\DP_OP_158_296_6262/n1176 ), 
	.B(\DP_OP_158_296_6262/n1198 ), 
	.A(\DP_OP_158_296_6262/n1178 ));
   NAND2X1TS U1725 (.Y(\DP_OP_158_296_6262/n1132 ), 
	.B(\DP_OP_158_296_6262/n1134 ), 
	.A(\DP_OP_158_296_6262/n1158 ));
   NAND2X1TS U1726 (.Y(\DP_OP_158_296_6262/n1075 ), 
	.B(\DP_OP_158_296_6262/n1109 ), 
	.A(\DP_OP_158_296_6262/n1077 ));
   NAND2X2TS U1727 (.Y(\DP_OP_158_296_6262/n912 ), 
	.B(n1471), 
	.A(\DP_OP_158_296_6262/n931 ));
   NOR2X4TS U1728 (.Y(\DP_OP_158_296_6262/n897 ), 
	.B(\DP_OP_158_296_6262/n899 ), 
	.A(\DP_OP_158_296_6262/n912 ));
   NAND2X6TS U1729 (.Y(\DP_OP_158_296_6262/n895 ), 
	.B(\DP_OP_158_296_6262/n956 ), 
	.A(\DP_OP_158_296_6262/n897 ));
   OR2X8TS U1730 (.Y(\addr_calc/fft_read_calc/counter/N38 ), 
	.B(\DP_OP_158_296_6262/n1071 ), 
	.A(\DP_OP_158_296_6262/n895 ));
   AOI21X4TS U1731 (.Y(n2794), 
	.B0(n2588), 
	.A1(FE_OFN333_data_to_fft), 
	.A0(\addr_calc/fft_read_calc/counter/N38 ));
   AOI2BB1X4TS U1733 (.Y(\addr_calc/iir_write_addr[27] ), 
	.B0(n1604), 
	.A1N(n1603), 
	.A0N(\add_x_19_5/n60 ));
   NAND2BX1TS U1734 (.Y(n1608), 
	.B(FE_OFN551_n1751), 
	.AN(n1609));
   NOR2X8TS U1735 (.Y(\DP_OP_158_296_6262/n1918 ), 
	.B(FE_OFN482_filesize_16_), 
	.A(FE_OFN480_filesize_17_));
   INVX6TS U1736 (.Y(n1611), 
	.A(\add_x_19_4/n69 ));
   OAI21X2TS U1738 (.Y(\add_x_19_4/n50 ), 
	.B0(\add_x_19_4/n52 ), 
	.A1(\add_x_19_4/n51 ), 
	.A0(FE_OCPN1230_n1611));
   OAI21X4TS U1739 (.Y(\add_x_19_4/n65 ), 
	.B0(\add_x_19_4/n67 ), 
	.A1(\add_x_19_4/n66 ), 
	.A0(FE_OCPN1230_n1611));
   NAND2X4TS U1740 (.Y(\DP_OP_158_296_6262/n1903 ), 
	.B(\DP_OP_158_296_6262/n1906 ), 
	.A(\DP_OP_158_296_6262/n1918 ));
   INVXLTS U1741 (.Y(\DP_OP_158_296_6262/n1891 ), 
	.A(\DP_OP_158_296_6262/n1890 ));
   XNOR2X4TS U1742 (.Y(n1730), 
	.B(FE_OFN473_filesize_23_), 
	.A(\DP_OP_158_296_6262/n1881 ));
   AOI21X4TS U1743 (.Y(n2805), 
	.B0(n2061), 
	.A1(FE_OFN319_data_from_fir), 
	.A0(\addr_calc/fir_write_calc/counter/N38 ));
   NAND2BXLTS U1744 (.Y(n1612), 
	.B(FE_OFN59_n2807), 
	.AN(n1613));
   NAND2X1TS U1745 (.Y(n1617), 
	.B(\addr_calc/fir_write_calc/counter/N73 ), 
	.A(FE_OFN549_n1763));
   OAI2BB1X1TS U1746 (.Y(n1100), 
	.B0(n1617), 
	.A1N(FE_OCPUNCON1090_n2805), 
	.A0N(FE_OFN238_addr_calc_fir_write_calc_count_30_));
   NAND2BX1TS U1747 (.Y(n1618), 
	.B(n1763), 
	.AN(n1619));
   OAI2BB1X1TS U1748 (.Y(n1023), 
	.B0(n1620), 
	.A1N(n2794), 
	.A0N(n1970));
   INVX2TS U1749 (.Y(\DP_OP_159_297_3515/n861 ), 
	.A(FE_OFN472_filesize_23_));
   NAND2X2TS U1750 (.Y(\DP_OP_159_297_3515/n941 ), 
	.B(\DP_OP_159_297_3515/n942 ), 
	.A(FE_OCPUNCON1565_n1789));
   XOR2X4TS U1751 (.Y(\DP_OP_159_297_3515/n1133 ), 
	.B(\DP_OP_159_297_3515/n861 ), 
	.A(\DP_OP_159_297_3515/n941 ));
   XOR2X2TS U1752 (.Y(\DP_OP_159_297_3515/n144 ), 
	.B(\add_x_22_4/n33 ), 
	.A(n1703));
   XOR2X4TS U1753 (.Y(\DP_OP_159_297_3515/n157 ), 
	.B(n1923), 
	.A(n1699));
   XNOR2X2TS U1755 (.Y(\DP_OP_159_297_3515/n70 ), 
	.B(FE_OFN235_addr_calc_iir_read_calc_count_27_), 
	.A(n1702));
   XOR2X4TS U1756 (.Y(\DP_OP_159_297_3515/n102 ), 
	.B(n1925), 
	.A(n1732));
   NOR2X2TS U1757 (.Y(\DP_OP_159_297_3515/n114 ), 
	.B(\DP_OP_159_297_3515/n116 ), 
	.A(\DP_OP_159_297_3515/n131 ));
   NOR2X4TS U1758 (.Y(\DP_OP_159_297_3515/n142 ), 
	.B(\DP_OP_159_297_3515/n157 ), 
	.A(\DP_OP_159_297_3515/n144 ));
   NOR2X2TS U1759 (.Y(\DP_OP_159_297_3515/n49 ), 
	.B(\DP_OP_159_297_3515/n51 ), 
	.A(\DP_OP_159_297_3515/n70 ));
   NAND2X2TS U1760 (.Y(\DP_OP_159_297_3515/n112 ), 
	.B(\DP_OP_159_297_3515/n142 ), 
	.A(\DP_OP_159_297_3515/n114 ));
   NAND2X4TS U1761 (.Y(\DP_OP_159_297_3515/n47 ), 
	.B(\DP_OP_159_297_3515/n49 ), 
	.A(\DP_OP_159_297_3515/n85 ));
   NOR2X6TS U1762 (.Y(\DP_OP_159_297_3515/n3 ), 
	.B(\DP_OP_159_297_3515/n5 ), 
	.A(\DP_OP_159_297_3515/n18 ));
   NOR2X4TS U1763 (.Y(\DP_OP_159_297_3515/n45 ), 
	.B(\DP_OP_159_297_3515/n112 ), 
	.A(\DP_OP_159_297_3515/n47 ));
   NAND2X4TS U1764 (.Y(\DP_OP_159_297_3515/n1 ), 
	.B(\DP_OP_159_297_3515/n3 ), 
	.A(\DP_OP_159_297_3515/n45 ));
   NOR2BX4TS U1765 (.Y(n2795), 
	.B(n1675), 
	.AN(n1625));
   OAI2BB1X1TS U1766 (.Y(n1013), 
	.B0(n1627), 
	.A1N(FE_OFN11_n2794), 
	.A0N(\addr_calc/fft_read_calc/count[21] ));
   NAND2BX1TS U1767 (.Y(n1630), 
	.B(FE_OFN3_n1754), 
	.AN(n1631));
   OAI2BB1X1TS U1768 (.Y(n1008), 
	.B0(n1630), 
	.A1N(FE_OFN12_n2794), 
	.A0N(n2575));
   INVX1TS U1769 (.Y(n1632), 
	.A(\add_x_19_4/n128 ));
   NAND2BX1TS U1770 (.Y(n1633), 
	.B(n1751), 
	.AN(n1634));
   OAI2BB1X1TS U1771 (.Y(n1017), 
	.B0(n1633), 
	.A1N(FE_OFN9_n2794), 
	.A0N(\addr_calc/fft_read_calc/count[17] ));
   NOR2X4TS U1772 (.Y(n1797), 
	.B(FE_OFN502_filesize_0_), 
	.A(FE_OFN501_filesize_1_));
   CLKINVX1TS U1774 (.Y(\add_x_19_4/n208 ), 
	.A(\add_x_19_4/n120 ));
   NAND2BX1TS U1775 (.Y(n1636), 
	.B(FE_OFN2_n1754), 
	.AN(n1637));
   OAI2BB1X1TS U1776 (.Y(n1016), 
	.B0(n1636), 
	.A1N(FE_OFN10_n2794), 
	.A0N(n2569));
   NAND2BX1TS U1777 (.Y(n1638), 
	.B(FE_OFN6_n1750), 
	.AN(n1639));
   OAI2BB1X1TS U1778 (.Y(n1018), 
	.B0(n1638), 
	.A1N(FE_OFN9_n2794), 
	.A0N(n2554));
   INVX2TS U1780 (.Y(\add_x_19_4/n40 ), 
	.A(\add_x_19_4/n42 ));
   INVX1TS U1782 (.Y(\add_x_19_4/n198 ), 
	.A(\add_x_19_4/n63 ));
   CLKINVX1TS U1783 (.Y(\add_x_19_4/n195 ), 
	.A(\add_x_19_4/n48 ));
   XOR2X2TS U1784 (.Y(\DP_OP_158_296_6262/n2056 ), 
	.B(n1664), 
	.A(\DP_OP_158_296_6262/n1860 ));
   XOR2X4TS U1785 (.Y(n1776), 
	.B(\DP_OP_158_296_6262/n1897 ), 
	.A(n1642));
   NAND2BX1TS U1786 (.Y(n1643), 
	.B(FE_OFN551_n1751), 
	.AN(n1644));
   OAI2BB1X2TS U1787 (.Y(n1030), 
	.B0(n1643), 
	.A1N(FE_OFN15_n2794), 
	.A0N(\addr_calc/fft_read_calc/count[4] ));
   NAND2BX1TS U1788 (.Y(n1645), 
	.B(FE_OFN69_n2809), 
	.AN(n1837));
   NAND2BX1TS U1789 (.Y(n1646), 
	.B(FE_OFN548_n1763), 
	.AN(n1647));
   OAI2BB1X1TS U1790 (.Y(n1118), 
	.B0(n1646), 
	.A1N(FE_OCPUNCON1084_n2805), 
	.A0N(FE_OFN233_addr_calc_fir_write_calc_count_12_));
   NOR2X2TS U1791 (.Y(\DP_OP_159_297_3515/n1075 ), 
	.B(FE_OFN499_filesize_2_), 
	.A(FE_OFN500_filesize_1_));
   NAND2X1TS U1792 (.Y(\DP_OP_159_297_3515/n1066 ), 
	.B(FE_OFN496_filesize_4_), 
	.A(FE_OFN498_filesize_3_));
   XOR2X2TS U1793 (.Y(n2607), 
	.B(\DP_OP_159_297_3515/n867 ), 
	.A(FE_OFN553_n1789));
   AO22X1TS U1795 (.Y(n985), 
	.B1(FE_OCPUNCON1570_n2812), 
	.B0(n1954), 
	.A1(\addr_calc/iir_write_calc/counter/N60 ), 
	.A0(FE_OCPUNCON1882_n2813));
   AO22X1TS U1797 (.Y(n979), 
	.B1(\addr_calc/iir_write_calc/count[23] ), 
	.B0(FE_OCPUNCON1572_n2812), 
	.A1(\addr_calc/iir_write_calc/counter/N66 ), 
	.A0(FE_OCPUNCON1884_n2813));
   AO22X1TS U1798 (.Y(n1136), 
	.B1(\addr_calc/iir_write_calc/count[31] ), 
	.B0(FE_OCPUNCON1575_n2812), 
	.A1(\addr_calc/iir_write_calc/counter/N74 ), 
	.A0(FE_OCPUNCON1886_n2813));
   AO22X1TS U1801 (.Y(n1001), 
	.B1(n1931), 
	.B0(FE_OCPUNCON1575_n2812), 
	.A1(\addr_calc/iir_write_calc/counter/N44 ), 
	.A0(FE_OCPUNCON1887_n2813));
   AO22X1TS U1802 (.Y(n978), 
	.B1(\addr_calc/iir_write_calc/count[24] ), 
	.B0(FE_OCPUNCON1573_n2812), 
	.A1(\addr_calc/iir_write_calc/counter/N67 ), 
	.A0(FE_OCPUNCON1886_n2813));
   AO22X1TS U1803 (.Y(n999), 
	.B1(\addr_calc/iir_write_calc/count[3] ), 
	.B0(FE_OCPUNCON1575_n2812), 
	.A1(\addr_calc/iir_write_calc/counter/N46 ), 
	.A0(FE_OCPUNCON1887_n2813));
   AO22X4TS U1804 (.Y(n997), 
	.B1(n1686), 
	.B0(FE_OCPUNCON1576_n2812), 
	.A1(\addr_calc/iir_write_calc/counter/N48 ), 
	.A0(FE_OCPUNCON1888_n2813));
   NOR2X2TS U1805 (.Y(n2813), 
	.B(n787), 
	.A(n1468));
   NOR2X2TS U1806 (.Y(n2790), 
	.B(n2788), 
	.A(n2789));
   INVX2TS U1807 (.Y(n1740), 
	.A(FE_OCPUNCON1570_n2812));
   OAI2BB2XLTS U1808 (.Y(n1000), 
	.B1(\add_x_22_5/n117 ), 
	.B0(n1740), 
	.A1N(\addr_calc/iir_write_calc/counter/N45 ), 
	.A0N(FE_OCPUNCON1887_n2813));
   NAND2X1TS U1809 (.Y(\DP_OP_159_297_3515/n927 ), 
	.B(\DP_OP_159_297_3515/n928 ), 
	.A(n1792));
   NAND2X2TS U1810 (.Y(\DP_OP_159_297_3515/n955 ), 
	.B(\DP_OP_159_297_3515/n956 ), 
	.A(n1792));
   XOR2X4TS U1813 (.Y(n1732), 
	.B(FE_OFN470_filesize_25_), 
	.A(\DP_OP_159_297_3515/n927 ));
   OAI2BB2XLTS U1814 (.Y(n974), 
	.B1(n1973), 
	.B0(n1740), 
	.A1N(\addr_calc/iir_write_calc/counter/N71 ), 
	.A0N(FE_OCPUNCON1884_n2813));
   NOR4X1TS U1815 (.Y(n796), 
	.D(n926), 
	.C(n925), 
	.B(iir_write_done), 
	.A(n1478));
   XNOR2X1TS U1818 (.Y(\DP_OP_158_296_6262/n174 ), 
	.B(n1985), 
	.A(n1776));
   XNOR2X4TS U1820 (.Y(n1651), 
	.B(n2362), 
	.A(\DP_OP_158_296_6262/n1991 ));
   XNOR2X4TS U1821 (.Y(n1654), 
	.B(FE_OFN478_filesize_19_), 
	.A(\DP_OP_158_296_6262/n1909 ));
   XNOR2X4TS U1822 (.Y(n1656), 
	.B(n2367), 
	.A(\DP_OP_158_296_6262/n1971 ));
   XNOR2X4TS U1823 (.Y(n1657), 
	.B(FE_OFN486_filesize_14_), 
	.A(\DP_OP_158_296_6262/n1943 ));
   XNOR2X4TS U1824 (.Y(n1658), 
	.B(FE_OFN484_filesize_15_), 
	.A(\DP_OP_158_296_6262/n1936 ));
   XNOR2X4TS U1825 (.Y(n1660), 
	.B(n1681), 
	.A(\DP_OP_158_296_6262/n1964 ));
   XNOR2X4TS U1826 (.Y(n1661), 
	.B(n2343), 
	.A(\DP_OP_159_297_3515/n920 ));
   AOI21X4TS U1827 (.Y(\add_x_19_4/n102 ), 
	.B0(\add_x_19_4/n104 ), 
	.A1(\add_x_19_4/n103 ), 
	.A0(\add_x_19_4/n112 ));
   NAND2X1TS U1830 (.Y(\DP_OP_159_297_3515/n1010 ), 
	.B(\DP_OP_159_297_3515/n1011 ), 
	.A(n1788));
   XNOR2X4TS U1831 (.Y(n2617), 
	.B(\DP_OP_159_297_3515/n870 ), 
	.A(\DP_OP_159_297_3515/n1003 ));
   CLKXOR2X2TS U1832 (.Y(\DP_OP_158_296_6262/n2034 ), 
	.B(n2371), 
	.A(\DP_OP_158_296_6262/n2010 ));
   NOR2X2TS U1833 (.Y(\DP_OP_158_296_6262/n1874 ), 
	.B(\DP_OP_158_296_6262/n1875 ), 
	.A(n1717));
   NAND2X2TS U1834 (.Y(\DP_OP_159_297_3515/n948 ), 
	.B(\DP_OP_159_297_3515/n949 ), 
	.A(n1792));
   INVX2TS U1839 (.Y(n1755), 
	.A(n1701));
   INVX4TS U1840 (.Y(\add_x_19_2/n91 ), 
	.A(\add_x_19_2/n92 ));
   CLKINVX2TS U1841 (.Y(\add_x_22_2/n23 ), 
	.A(\add_x_22_2/n24 ));
   CLKINVX2TS U1842 (.Y(\add_x_22_5/n23 ), 
	.A(\add_x_22_5/n24 ));
   CLKINVX2TS U1843 (.Y(\add_x_22_3/n23 ), 
	.A(\add_x_22_3/n24 ));
   CLKINVX2TS U1844 (.Y(\add_x_22_5/n75 ), 
	.A(\add_x_22_5/n76 ));
   INVX2TS U1845 (.Y(\add_x_22_4/n23 ), 
	.A(\add_x_22_4/n24 ));
   CLKINVX2TS U1846 (.Y(\add_x_22_4/n41 ), 
	.A(\add_x_22_4/n42 ));
   CLKINVX2TS U1847 (.Y(\add_x_22_3/n75 ), 
	.A(\add_x_22_3/n76 ));
   INVX1TS U1848 (.Y(\add_x_22_4/n75 ), 
	.A(\add_x_22_4/n76 ));
   CLKINVX2TS U1849 (.Y(\add_x_22_1/n23 ), 
	.A(\add_x_22_1/n24 ));
   XNOR2X1TS U1850 (.Y(\DP_OP_158_296_6262/n277 ), 
	.B(n1994), 
	.A(n1756));
   INVX2TS U1851 (.Y(\add_x_22_0/n93 ), 
	.A(\add_x_22_0/n94 ));
   NOR2X2TS U1852 (.Y(\add_x_19_4/n72 ), 
	.B(\add_x_19_4/n93 ), 
	.A(\add_x_19_4/n74 ));
   CLKINVX2TS U1853 (.Y(\add_x_19_3/n177 ), 
	.A(\add_x_19_3/n178 ));
   NOR2X1TS U1854 (.Y(\DP_OP_159_297_3515/n921 ), 
	.B(n1155), 
	.A(\DP_OP_159_297_3515/n852 ));
   CLKINVX1TS U1855 (.Y(\add_x_22_5/n118 ), 
	.A(\add_x_22_5/n119 ));
   INVX1TS U1856 (.Y(\add_x_19_3/n174 ), 
	.A(\add_x_19_3/n176 ));
   CLKINVX1TS U1857 (.Y(\add_x_19_4/n143 ), 
	.A(\add_x_19_4/n145 ));
   INVX1TS U1858 (.Y(\DP_OP_159_297_3515/n862 ), 
	.A(FE_OFN474_filesize_22_));
   INVX1TS U1859 (.Y(\add_x_19_1/n213 ), 
	.A(\add_x_19_1/n144 ));
   CLKINVX1TS U1860 (.Y(\add_x_19_1/n143 ), 
	.A(\add_x_19_1/n145 ));
   CLKINVX1TS U1861 (.Y(\add_x_19_0/n219 ), 
	.A(\add_x_19_0/n175 ));
   CLKINVX1TS U1862 (.Y(\add_x_19_3/n195 ), 
	.A(\add_x_19_3/n48 ));
   CLKINVX1TS U1863 (.Y(\add_x_19_1/n195 ), 
	.A(\add_x_19_1/n48 ));
   INVX1TS U1864 (.Y(\add_x_19_0/n195 ), 
	.A(\add_x_19_0/n48 ));
   INVX2TS U1866 (.Y(n1902), 
	.A(n1901));
   INVX2TS U1867 (.Y(n2046), 
	.A(n2045));
   INVX4TS U1868 (.Y(n1666), 
	.A(n1975));
   INVX2TS U1869 (.Y(n1907), 
	.A(\addr_calc/iir_read_calc/count[9] ));
   INVX2TS U1870 (.Y(n2024), 
	.A(\addr_calc/iir_read_calc/count[18] ));
   INVX2TS U1872 (.Y(\add_x_22_5/n67 ), 
	.A(\addr_calc/iir_write_calc/count[14] ));
   INVX2TS U1874 (.Y(n1921), 
	.A(\addr_calc/fft_write_calc/count[19] ));
   INVX2TS U1875 (.Y(n1891), 
	.A(\addr_calc/fir_write_calc/count[21] ));
   INVX2TS U1876 (.Y(n1981), 
	.A(\addr_calc/fir_read_calc/count[22] ));
   INVX2TS U1877 (.Y(n1938), 
	.A(\addr_calc/iir_write_calc/count[7] ));
   CLKINVX6TS U1891 (.Y(\add_x_19_3/n68 ), 
	.A(\add_x_19_3/n69 ));
   NAND2X1TS U1892 (.Y(n1735), 
	.B(n1681), 
	.A(n1733));
   INVX1TS U1893 (.Y(\add_x_22_2/n75 ), 
	.A(\add_x_22_2/n76 ));
   INVX1TS U1894 (.Y(\add_x_22_0/n75 ), 
	.A(\add_x_22_0/n76 ));
   INVX1TS U1895 (.Y(\add_x_22_1/n75 ), 
	.A(\add_x_22_1/n76 ));
   NOR2X4TS U1897 (.Y(\add_x_19_3/n46 ), 
	.B(\add_x_19_3/n48 ), 
	.A(\add_x_19_3/n51 ));
   INVX3TS U1900 (.Y(\add_x_19_0/n177 ), 
	.A(\add_x_19_0/n178 ));
   NAND2X4TS U1901 (.Y(\add_x_19_3/n51 ), 
	.B(\add_x_19_3/n53 ), 
	.A(\add_x_19_3/n61 ));
   INVX1TS U1904 (.Y(\add_x_19_2/n148 ), 
	.A(\add_x_19_2/n150 ));
   INVX1TS U1905 (.Y(\add_x_19_1/n148 ), 
	.A(\add_x_19_1/n150 ));
   INVX1TS U1906 (.Y(\add_x_19_3/n148 ), 
	.A(\add_x_19_3/n150 ));
   INVX1TS U1907 (.Y(\add_x_19_0/n148 ), 
	.A(\add_x_19_0/n150 ));
   INVX1TS U1908 (.Y(\add_x_19_2/n177 ), 
	.A(\add_x_19_2/n178 ));
   INVX1TS U1909 (.Y(\add_x_19_0/n186 ), 
	.A(\add_x_19_0/n187 ));
   INVX1TS U1910 (.Y(\add_x_19_5/n195 ), 
	.A(\add_x_19_5/n48 ));
   CLKINVX1TS U1911 (.Y(\add_x_19_4/n196 ), 
	.A(\add_x_19_4/n55 ));
   INVX2TS U1912 (.Y(n2061), 
	.A(FE_OFN566_n2066));
   INVX1TS U1914 (.Y(\add_x_19_2/n109 ), 
	.A(\add_x_19_2/n111 ));
   INVX1TS U1915 (.Y(\add_x_19_2/n186 ), 
	.A(\add_x_19_2/n187 ));
   INVX1TS U1916 (.Y(\add_x_19_2/n213 ), 
	.A(\add_x_19_2/n144 ));
   INVX1TS U1917 (.Y(\add_x_19_3/n186 ), 
	.A(\add_x_19_3/n187 ));
   NOR2X4TS U1918 (.Y(\add_x_19_0/n53 ), 
	.B(\add_x_19_0/n55 ), 
	.A(\add_x_19_0/n58 ));
   NOR2X2TS U1919 (.Y(\add_x_19_4/n151 ), 
	.B(FE_OFN424_offset_9_), 
	.A(n1685));
   INVX1TS U1920 (.Y(\add_x_19_5/n186 ), 
	.A(FE_OCPN1907_add_x_19_5_n187));
   INVX1TS U1921 (.Y(\add_x_19_5/n219 ), 
	.A(\add_x_19_5/n175 ));
   INVX1TS U1922 (.Y(\add_x_19_1/n109 ), 
	.A(\add_x_19_1/n111 ));
   NOR2X1TS U1923 (.Y(\add_x_19_4/n76 ), 
	.B(\add_x_19_4/n81 ), 
	.A(\add_x_19_4/n78 ));
   NOR2X2TS U1924 (.Y(\add_x_19_5/n103 ), 
	.B(\add_x_19_5/n105 ), 
	.A(\add_x_19_5/n110 ));
   INVX1TS U1925 (.Y(\add_x_19_4/n222 ), 
	.A(\add_x_19_4/n188 ));
   INVX1TS U1926 (.Y(\add_x_19_5/n222 ), 
	.A(\add_x_19_5/n188 ));
   INVX1TS U1927 (.Y(\add_x_19_0/n213 ), 
	.A(\add_x_19_0/n144 ));
   INVX1TS U1928 (.Y(\add_x_19_1/n219 ), 
	.A(\add_x_19_1/n175 ));
   INVX1TS U1929 (.Y(\add_x_19_0/n109 ), 
	.A(\add_x_19_0/n111 ));
   INVX1TS U1930 (.Y(\add_x_19_4/n219 ), 
	.A(\add_x_19_4/n175 ));
   INVX2TS U1931 (.Y(n2365), 
	.A(\DP_OP_159_297_3515/n875 ));
   INVX2TS U1933 (.Y(n2364), 
	.A(\DP_OP_159_297_3515/n876 ));
   INVX2TS U1935 (.Y(n2366), 
	.A(\DP_OP_159_297_3515/n878 ));
   INVX2TS U1936 (.Y(n1838), 
	.A(n1837));
   INVX2TS U1938 (.Y(n1784), 
	.A(\add_x_22_4/n67 ));
   INVX2TS U1939 (.Y(n1983), 
	.A(n1982));
   INVX3TS U1940 (.Y(n1985), 
	.A(n1984));
   INVX2TS U1941 (.Y(n1690), 
	.A(n1991));
   INVX2TS U1942 (.Y(n2566), 
	.A(\add_x_22_4/n64 ));
   INVX2TS U1943 (.Y(n1835), 
	.A(n1834));
   INVX6TS U1944 (.Y(n1686), 
	.A(n1937));
   INVX2TS U1946 (.Y(n2043), 
	.A(n2042));
   INVX2TS U1947 (.Y(n1689), 
	.A(n1963));
   INVX1TS U1948 (.Y(\add_x_22_4/n109 ), 
	.A(\addr_calc/iir_read_calc/count[4] ));
   CLKINVX2TS U1949 (.Y(n1956), 
	.A(n1955));
   INVX2TS U1950 (.Y(n2569), 
	.A(\add_x_22_0/n49 ));
   INVX2TS U1951 (.Y(n1851), 
	.A(n1850));
   CLKINVX3TS U1952 (.Y(n2028), 
	.A(n2027));
   INVX2TS U1953 (.Y(n1664), 
	.A(n2343));
   NOR2X1TS U1954 (.Y(\DP_OP_158_296_6262/n1837 ), 
	.B(FE_OFN466_filesize_28_), 
	.A(FE_OFN465_filesize_29_));
   INVX2TS U1956 (.Y(\add_x_22_0/n114 ), 
	.A(\addr_calc/fft_read_calc/count[3] ));
   INVX2TS U1959 (.Y(n1937), 
	.A(\addr_calc/iir_write_calc/count[5] ));
   INVX2TS U1961 (.Y(n2047), 
	.A(\addr_calc/iir_write_calc/count[20] ));
   INVX2TS U1962 (.Y(n1665), 
	.A(n2040));
   INVX2TS U1964 (.Y(n1923), 
	.A(\addr_calc/iir_read_calc/count[21] ));
   INVX2TS U1965 (.Y(n1971), 
	.A(\addr_calc/iir_write_calc/count[27] ));
   INVX2TS U1967 (.Y(\add_x_22_0/n15 ), 
	.A(\addr_calc/fft_read_calc/count[26] ));
   INVX2TS U1969 (.Y(\add_x_22_4/n46 ), 
	.A(\addr_calc/iir_read_calc/count[19] ));
   INVX2TS U1970 (.Y(n1668), 
	.A(n2012));
   INVX2TS U1971 (.Y(n1984), 
	.A(\addr_calc/fir_read_calc/count[20] ));
   INVX2TS U1972 (.Y(n1899), 
	.A(\addr_calc/fir_read_calc/count[9] ));
   INVX2TS U1973 (.Y(n1870), 
	.A(\addr_calc/fir_read_calc/count[28] ));
   INVX2TS U1975 (.Y(n1841), 
	.A(\addr_calc/fir_read_calc/count[29] ));
   INVX2TS U1976 (.Y(n1837), 
	.A(\addr_calc/fir_read_calc/count[30] ));
   INVX4TS U2016 (.Y(n1763), 
	.A(n1758));
   CLKINVX3TS U2022 (.Y(n1675), 
	.A(\addr_calc/fft_write_calc/counter/N38 ));
   XNOR2X4TS U2024 (.Y(\addr_calc/fir_write_addr[28] ), 
	.B(\add_x_19_3/n4 ), 
	.A(\add_x_19_3/n50 ));
   OR3X1TS U2025 (.Y(n1696), 
	.C(FE_OFN562_n2060), 
	.B(n2808), 
	.A(FE_OFN329_data_cntl_N99));
   INVX2TS U2028 (.Y(\add_x_19_5/n133 ), 
	.A(\add_x_19_5/n134 ));
   INVX2TS U2029 (.Y(\add_x_19_1/n133 ), 
	.A(\add_x_19_1/n134 ));
   INVX3TS U2030 (.Y(\add_x_19_2/n133 ), 
	.A(\add_x_19_2/n134 ));
   INVX2TS U2031 (.Y(\add_x_19_3/n133 ), 
	.A(\add_x_19_3/n134 ));
   CLKINVX2TS U2032 (.Y(\add_x_22_0/n41 ), 
	.A(\add_x_22_0/n42 ));
   CLKINVX2TS U2033 (.Y(\add_x_22_1/n41 ), 
	.A(\add_x_22_1/n42 ));
   CLKINVX2TS U2034 (.Y(\add_x_22_2/n41 ), 
	.A(\add_x_22_2/n42 ));
   CLKINVX2TS U2035 (.Y(\add_x_22_3/n41 ), 
	.A(\add_x_22_3/n42 ));
   CLKINVX2TS U2036 (.Y(\add_x_22_5/n41 ), 
	.A(\add_x_22_5/n42 ));
   INVX1TS U2039 (.Y(\add_x_22_1/n58 ), 
	.A(\add_x_22_1/n59 ));
   INVX1TS U2040 (.Y(\add_x_22_4/n58 ), 
	.A(FE_OFN150_add_x_22_4_n59));
   INVX1TS U2041 (.Y(\add_x_22_5/n58 ), 
	.A(FE_OFN148_add_x_22_5_n59));
   OAI21X1TS U2042 (.Y(n2798), 
	.B0(n2073), 
	.A1(n2796), 
	.A0(\addr_calc/fft_write_calc/counter/N43 ));
   INVX1TS U2043 (.Y(\add_x_22_3/n58 ), 
	.A(\add_x_22_3/n59 ));
   INVX1TS U2044 (.Y(\add_x_22_0/n58 ), 
	.A(\add_x_22_0/n59 ));
   INVX1TS U2046 (.Y(\add_x_22_2/n58 ), 
	.A(FE_OFN147_add_x_22_2_n59));
   AOI21X4TS U2047 (.Y(\add_x_19_3/n52 ), 
	.B0(\add_x_19_3/n54 ), 
	.A1(\add_x_19_3/n53 ), 
	.A0(\add_x_19_3/n62 ));
   INVX2TS U2048 (.Y(n1830), 
	.A(n936));
   NAND2X1TS U2050 (.Y(\DP_OP_159_297_3515/n1031 ), 
	.B(n2365), 
	.A(n1787));
   CLKINVX2TS U2051 (.Y(\add_x_22_3/n93 ), 
	.A(\add_x_22_3/n94 ));
   CLKINVX2TS U2052 (.Y(\add_x_22_4/n93 ), 
	.A(\add_x_22_4/n94 ));
   CLKINVX2TS U2053 (.Y(\add_x_22_2/n93 ), 
	.A(\add_x_22_2/n94 ));
   OAI21X4TS U2054 (.Y(\add_x_19_3/n73 ), 
	.B0(\add_x_19_3/n75 ), 
	.A1(\add_x_19_3/n74 ), 
	.A0(\add_x_19_3/n94 ));
   CLKINVX2TS U2055 (.Y(\add_x_22_5/n93 ), 
	.A(FE_OFN149_add_x_22_5_n94));
   OAI21X1TS U2056 (.Y(n2792), 
	.B0(n2815), 
	.A1(n2790), 
	.A0(n2791));
   CLKINVX2TS U2057 (.Y(\add_x_22_1/n93 ), 
	.A(\add_x_22_1/n94 ));
   CLKINVX1TS U2058 (.Y(\add_x_19_0/n147 ), 
	.A(\add_x_19_0/n149 ));
   CLKINVX1TS U2059 (.Y(\add_x_19_1/n147 ), 
	.A(\add_x_19_1/n149 ));
   CLKINVX1TS U2060 (.Y(\add_x_19_2/n147 ), 
	.A(\add_x_19_2/n149 ));
   CLKINVX1TS U2061 (.Y(\add_x_19_3/n147 ), 
	.A(\add_x_19_3/n149 ));
   CLKINVX1TS U2062 (.Y(\add_x_19_5/n147 ), 
	.A(\add_x_19_5/n149 ));
   INVX1TS U2063 (.Y(\add_x_19_5/n148 ), 
	.A(\add_x_19_5/n150 ));
   INVX1TS U2064 (.Y(\add_x_19_4/n148 ), 
	.A(\add_x_19_4/n150 ));
   CLKINVX1TS U2065 (.Y(\add_x_19_4/n147 ), 
	.A(\add_x_19_4/n149 ));
   INVX1TS U2067 (.Y(\add_x_22_5/n110 ), 
	.A(\add_x_22_5/n111 ));
   INVX1TS U2068 (.Y(\add_x_22_3/n110 ), 
	.A(\add_x_22_3/n111 ));
   AOI21X4TS U2069 (.Y(\add_x_19_1/n94 ), 
	.B0(\add_x_19_1/n96 ), 
	.A1(\add_x_19_1/n95 ), 
	.A0(\add_x_19_1/n104 ));
   INVX2TS U2071 (.Y(\add_x_19_1/n177 ), 
	.A(\add_x_19_1/n178 ));
   AOI21X2TS U2073 (.Y(\add_x_19_0/n52 ), 
	.B0(\add_x_19_0/n54 ), 
	.A1(\add_x_19_0/n62 ), 
	.A0(\add_x_19_0/n53 ));
   INVX1TS U2074 (.Y(\add_x_22_0/n110 ), 
	.A(\add_x_22_0/n111 ));
   INVX1TS U2075 (.Y(\add_x_22_4/n110 ), 
	.A(\add_x_22_4/n111 ));
   CLKINVX1TS U2076 (.Y(\add_x_19_5/n214 ), 
	.A(\add_x_19_5/n151 ));
   INVX1TS U2077 (.Y(\DP_OP_159_297_3515/n928 ), 
	.A(\DP_OP_159_297_3515/n852 ));
   OAI21X2TS U2078 (.Y(\add_x_19_1/n150 ), 
	.B0(\add_x_19_1/n152 ), 
	.A1(\add_x_19_1/n155 ), 
	.A0(\add_x_19_1/n151 ));
   CLKINVX1TS U2079 (.Y(\add_x_19_0/n208 ), 
	.A(\add_x_19_0/n120 ));
   CLKINVX1TS U2080 (.Y(\add_x_19_0/n204 ), 
	.A(\add_x_19_0/n97 ));
   CLKINVX2TS U2081 (.Y(n2585), 
	.A(n2074));
   CLKINVX1TS U2082 (.Y(\add_x_19_3/n204 ), 
	.A(\add_x_19_3/n97 ));
   CLKINVX1TS U2083 (.Y(\add_x_19_4/n202 ), 
	.A(\add_x_19_4/n86 ));
   OAI21X4TS U2084 (.Y(\add_x_19_3/n104 ), 
	.B0(\add_x_19_3/n106 ), 
	.A1(\add_x_19_3/n111 ), 
	.A0(\add_x_19_3/n105 ));
   INVX1TS U2085 (.Y(\add_x_19_3/n208 ), 
	.A(\add_x_19_3/n120 ));
   CLKINVX1TS U2086 (.Y(\add_x_19_1/n202 ), 
	.A(\add_x_19_1/n86 ));
   CLKINVX1TS U2087 (.Y(\add_x_19_0/n202 ), 
	.A(\add_x_19_0/n86 ));
   CLKINVX1TS U2088 (.Y(\add_x_19_0/n210 ), 
	.A(\add_x_19_0/n128 ));
   CLKINVX1TS U2089 (.Y(\add_x_19_4/n206 ), 
	.A(\add_x_19_4/n105 ));
   CLKINVX1TS U2090 (.Y(\add_x_19_5/n202 ), 
	.A(\add_x_19_5/n86 ));
   INVX1TS U2091 (.Y(\add_x_19_4/n207 ), 
	.A(\add_x_19_4/n110 ));
   INVX1TS U2092 (.Y(\add_x_19_4/n109 ), 
	.A(\add_x_19_4/n111 ));
   INVX1TS U2093 (.Y(\add_x_22_0/n118 ), 
	.A(\add_x_22_0/n119 ));
   CLKINVX1TS U2094 (.Y(\add_x_19_3/n202 ), 
	.A(\add_x_19_3/n86 ));
   INVX1TS U2095 (.Y(\add_x_19_2/n207 ), 
	.A(\add_x_19_2/n110 ));
   INVX1TS U2096 (.Y(\add_x_22_4/n118 ), 
	.A(\add_x_22_4/n119 ));
   INVX1TS U2097 (.Y(\add_x_22_2/n110 ), 
	.A(\add_x_22_2/n111 ));
   CLKINVX1TS U2098 (.Y(\add_x_19_1/n198 ), 
	.A(\add_x_19_1/n63 ));
   INVX1TS U2099 (.Y(\add_x_22_1/n110 ), 
	.A(\add_x_22_1/n111 ));
   CLKINVX1TS U2100 (.Y(\add_x_19_4/n199 ), 
	.A(\add_x_19_4/n66 ));
   CLKINVX1TS U2101 (.Y(\add_x_19_3/n221 ), 
	.A(\add_x_19_3/n184 ));
   CLKINVX1TS U2102 (.Y(\add_x_19_0/n198 ), 
	.A(\add_x_19_0/n63 ));
   CLKINVX1TS U2103 (.Y(\add_x_19_5/n198 ), 
	.A(\add_x_19_5/n63 ));
   INVX1TS U2105 (.Y(\add_x_19_4/n186 ), 
	.A(\add_x_19_4/n187 ));
   NOR2X4TS U2107 (.Y(\add_x_19_2/n151 ), 
	.B(FE_OCPUNCON654_FE_OFN422_offset_9_), 
	.A(n1900));
   CLKAND2X2TS U2108 (.Y(n2603), 
	.B(n2341), 
	.A(FE_OFN465_filesize_29_));
   CLKINVX1TS U2109 (.Y(\add_x_19_5/n220 ), 
	.A(\add_x_19_5/n181 ));
   INVX1TS U2110 (.Y(\add_x_19_3/n219 ), 
	.A(\add_x_19_3/n175 ));
   CLKINVX1TS U2111 (.Y(\add_x_19_3/n217 ), 
	.A(\add_x_19_3/n165 ));
   INVX2TS U2112 (.Y(n1976), 
	.A(\add_x_22_1/n64 ));
   INVX1TS U2113 (.Y(\add_x_22_2/n118 ), 
	.A(\add_x_22_2/n119 ));
   INVX1TS U2114 (.Y(\add_x_22_3/n118 ), 
	.A(\add_x_22_3/n119 ));
   CLKINVX1TS U2115 (.Y(\add_x_19_4/n212 ), 
	.A(\add_x_19_4/n139 ));
   INVX1TS U2116 (.Y(\add_x_19_4/n213 ), 
	.A(\add_x_19_4/n144 ));
   INVX1TS U2117 (.Y(\add_x_22_1/n118 ), 
	.A(\add_x_22_1/n119 ));
   CLKINVX1TS U2118 (.Y(\add_x_19_1/n208 ), 
	.A(\add_x_19_1/n120 ));
   CLKINVX1TS U2119 (.Y(\add_x_19_3/n215 ), 
	.A(\add_x_19_3/n154 ));
   CLKINVX2TS U2120 (.Y(n2372), 
	.A(\DP_OP_159_297_3515/n815 ));
   NOR2X2TS U2121 (.Y(\add_x_19_1/n103 ), 
	.B(\add_x_19_1/n105 ), 
	.A(\add_x_19_1/n110 ));
   OAI21X4TS U2122 (.Y(\add_x_19_1/n104 ), 
	.B0(\add_x_19_1/n106 ), 
	.A1(\add_x_19_1/n105 ), 
	.A0(\add_x_19_1/n111 ));
   NOR2X2TS U2123 (.Y(\add_x_19_2/n53 ), 
	.B(\add_x_19_2/n55 ), 
	.A(\add_x_19_2/n58 ));
   OAI21X4TS U2124 (.Y(\add_x_19_4/n187 ), 
	.B0(\add_x_19_4/n189 ), 
	.A1(\add_x_19_4/n191 ), 
	.A0(\add_x_19_4/n188 ));
   INVX2TS U2125 (.Y(n2362), 
	.A(\DP_OP_159_297_3515/n877 ));
   INVX1TS U2126 (.Y(\add_x_19_5/n213 ), 
	.A(\add_x_19_5/n144 ));
   CLKINVX1TS U2127 (.Y(\add_x_19_4/n221 ), 
	.A(\add_x_19_4/n184 ));
   INVX1TS U2128 (.Y(\add_x_19_3/n213 ), 
	.A(\add_x_19_3/n144 ));
   CLKINVX1TS U2129 (.Y(\add_x_19_2/n212 ), 
	.A(\add_x_19_2/n139 ));
   CLKINVX1TS U2130 (.Y(\DP_OP_159_297_3515/n944 ), 
	.A(\DP_OP_159_297_3515/n943 ));
   CLKINVX1TS U2131 (.Y(\add_x_19_5/n210 ), 
	.A(\add_x_19_5/n128 ));
   CLKINVX2TS U2132 (.Y(n1678), 
	.A(FE_OFN467_filesize_27_));
   CLKINVX1TS U2133 (.Y(\add_x_19_1/n174 ), 
	.A(\add_x_19_1/n176 ));
   CLKINVX1TS U2134 (.Y(\DP_OP_159_297_3515/n1025 ), 
	.A(\DP_OP_159_297_3515/n1026 ));
   CLKINVX1TS U2135 (.Y(\add_x_19_3/n218 ), 
	.A(\add_x_19_3/n170 ));
   CLKINVX1TS U2136 (.Y(\add_x_19_4/n217 ), 
	.A(\add_x_19_4/n165 ));
   INVX2TS U2137 (.Y(n2369), 
	.A(\DP_OP_159_297_3515/n867 ));
   CLKINVX1TS U2138 (.Y(\add_x_19_2/n215 ), 
	.A(\add_x_19_2/n154 ));
   CLKINVX1TS U2139 (.Y(\add_x_19_0/n215 ), 
	.A(\add_x_19_0/n154 ));
   CLKINVX1TS U2140 (.Y(\add_x_19_2/n210 ), 
	.A(\add_x_19_2/n128 ));
   INVX1TS U2141 (.Y(\add_x_19_2/n219 ), 
	.A(\add_x_19_2/n175 ));
   CLKINVX1TS U2142 (.Y(\add_x_19_2/n208 ), 
	.A(\add_x_19_2/n120 ));
   INVX1TS U2143 (.Y(\add_x_19_3/n207 ), 
	.A(\add_x_19_3/n110 ));
   INVX1TS U2144 (.Y(\add_x_19_0/n207 ), 
	.A(\add_x_19_0/n110 ));
   INVX1TS U2145 (.Y(\add_x_19_3/n198 ), 
	.A(\add_x_19_3/n63 ));
   CLKINVX1TS U2146 (.Y(\add_x_19_5/n206 ), 
	.A(\add_x_19_5/n105 ));
   CLKINVX1TS U2147 (.Y(\add_x_19_2/n206 ), 
	.A(\add_x_19_2/n105 ));
   INVX1TS U2148 (.Y(\add_x_19_5/n207 ), 
	.A(\add_x_19_5/n110 ));
   CLKINVX2TS U2149 (.Y(\add_x_19_5/n109 ), 
	.A(\add_x_19_5/n111 ));
   CLKINVX1TS U2150 (.Y(\add_x_19_1/n210 ), 
	.A(\add_x_19_1/n128 ));
   CLKINVX1TS U2151 (.Y(\add_x_19_2/n204 ), 
	.A(\add_x_19_2/n97 ));
   CLKINVX1TS U2152 (.Y(\add_x_19_1/n207 ), 
	.A(\add_x_19_1/n110 ));
   CLKINVX1TS U2153 (.Y(\add_x_19_4/n204 ), 
	.A(\add_x_19_4/n97 ));
   INVX2TS U2155 (.Y(n1990), 
	.A(n1989));
   INVX2TS U2156 (.Y(n2025), 
	.A(n2024));
   INVX2TS U2157 (.Y(n1895), 
	.A(\add_x_22_2/n80 ));
   INVX2TS U2158 (.Y(n1994), 
	.A(\add_x_22_2/n74 ));
   CLKINVX1TS U2159 (.Y(n2072), 
	.A(FE_OFN567_n2070));
   INVX2TS U2160 (.Y(n1880), 
	.A(\add_x_22_3/n71 ));
   INVX4TS U2161 (.Y(fir_enable), 
	.A(n2065));
   INVX2TS U2162 (.Y(n2007), 
	.A(n2810));
   INVX2TS U2163 (.Y(n1874), 
	.A(\add_x_22_3/n84 ));
   INVX2TS U2164 (.Y(n1883), 
	.A(n1882));
   INVX2TS U2165 (.Y(n1867), 
	.A(\add_x_22_3/n105 ));
   INVX2TS U2166 (.Y(n1872), 
	.A(\add_x_22_3/n89 ));
   INVX2TS U2167 (.Y(n1869), 
	.A(\add_x_22_3/n98 ));
   INVX2TS U2168 (.Y(n1866), 
	.A(\add_x_22_3/n114 ));
   INVX2TS U2169 (.Y(n1916), 
	.A(\add_x_22_4/n57 ));
   INVX2TS U2170 (.Y(n2074), 
	.A(FE_OFN567_n2070));
   INVX3TS U2171 (.Y(n1920), 
	.A(n1919));
   INVX2TS U2172 (.Y(n2041), 
	.A(\add_x_22_5/n92 ));
   INVX2TS U2173 (.Y(n1997), 
	.A(\add_x_22_2/n92 ));
   INVX2TS U2174 (.Y(n1908), 
	.A(\add_x_22_2/n114 ));
   INVX2TS U2176 (.Y(n1935), 
	.A(\add_x_22_5/n109 ));
   INVX2TS U2177 (.Y(n1945), 
	.A(\add_x_22_5/n71 ));
   INVX2TS U2179 (.Y(n1951), 
	.A(\add_x_22_5/n57 ));
   INVX2TS U2180 (.Y(n1879), 
	.A(n1878));
   INVX2TS U2181 (.Y(n1954), 
	.A(\add_x_22_5/n53 ));
   INVX2TS U2182 (.Y(n1888), 
	.A(n1887));
   INVX2TS U2183 (.Y(n1906), 
	.A(\add_x_22_2/n109 ));
   INVX2TS U2184 (.Y(n2020), 
	.A(n2019));
   INVX2TS U2185 (.Y(n2001), 
	.A(\add_x_22_2/n101 ));
   INVX2TS U2186 (.Y(n2044), 
	.A(\add_x_22_5/n74 ));
   INVX2TS U2187 (.Y(n1942), 
	.A(\add_x_22_5/n80 ));
   INVX2TS U2188 (.Y(n1896), 
	.A(\add_x_22_3/n7 ));
   INVX2TS U2190 (.Y(n1940), 
	.A(\add_x_22_5/n84 ));
   INVX2TS U2192 (.Y(n1842), 
	.A(n1841));
   INVX2TS U2193 (.Y(n1881), 
	.A(\add_x_22_2/n46 ));
   INVX2TS U2194 (.Y(n1884), 
	.A(\add_x_22_2/n53 ));
   INVX2TS U2195 (.Y(n1893), 
	.A(\add_x_22_2/n71 ));
   INVX2TS U2196 (.Y(n2039), 
	.A(\add_x_22_5/n101 ));
   INVX2TS U2197 (.Y(n1890), 
	.A(\add_x_22_2/n64 ));
   INVX2TS U2198 (.Y(n1932), 
	.A(\add_x_22_1/n84 ));
   INVX2TS U2199 (.Y(\add_x_22_1/n64 ), 
	.A(\addr_calc/fft_write_calc/count[15] ));
   CLKINVX1TS U2200 (.Y(\addr_calc/fft_write_calc/counter/N43 ), 
	.A(\addr_calc/fft_write_calc/count[0] ));
   INVX2TS U2201 (.Y(n1927), 
	.A(\add_x_22_1/n71 ));
   INVX1TS U2202 (.Y(\add_x_22_4/n84 ), 
	.A(\addr_calc/iir_read_calc/count[10] ));
   CLKINVX1TS U2203 (.Y(\add_x_22_4/n98 ), 
	.A(\addr_calc/iir_read_calc/count[7] ));
   INVX2TS U2204 (.Y(n2023), 
	.A(\add_x_22_1/n74 ));
   INVX2TS U2206 (.Y(n2049), 
	.A(\add_x_22_0/n92 ));
   INVX2TS U2208 (.Y(n2063), 
	.A(n2062));
   CLKINVX1TS U2209 (.Y(\add_x_22_4/n80 ), 
	.A(\addr_calc/iir_read_calc/count[11] ));
   INVX2TS U2210 (.Y(n1829), 
	.A(n1828));
   CLKINVX1TS U2211 (.Y(\add_x_22_1/n67 ), 
	.A(FE_OFN258_addr_calc_fft_write_calc_count_14_));
   INVX2TS U2212 (.Y(n1853), 
	.A(n1852));
   INVX1TS U2213 (.Y(\add_x_22_0/n109 ), 
	.A(FE_OFN263_addr_calc_fft_read_calc_count_4_));
   CLKINVX1TS U2214 (.Y(\add_x_22_0/n105 ), 
	.A(\addr_calc/fft_read_calc/count[5] ));
   INVX3TS U2215 (.Y(n2058), 
	.A(n2057));
   CLKINVX1TS U2217 (.Y(\add_x_22_3/n101 ), 
	.A(\addr_calc/fir_write_calc/count[6] ));
   INVX1TS U2218 (.Y(\add_x_22_3/n109 ), 
	.A(\addr_calc/fir_write_calc/count[4] ));
   INVX1TS U2219 (.Y(n1944), 
	.A(n1943));
   CLKINVX1TS U2220 (.Y(\add_x_22_3/n92 ), 
	.A(FE_OFN256_addr_calc_fir_write_calc_count_8_));
   INVX2TS U2221 (.Y(n2031), 
	.A(\add_x_22_4/n33 ));
   INVX2TS U2222 (.Y(n1936), 
	.A(\add_x_22_1/n98 ));
   INVX2TS U2224 (.Y(n2026), 
	.A(\add_x_22_1/n92 ));
   INVX2TS U2225 (.Y(n1934), 
	.A(\add_x_22_1/n89 ));
   INVX2TS U2226 (.Y(n2018), 
	.A(\add_x_22_4/n101 ));
   INVX2TS U2227 (.Y(n1924), 
	.A(\add_x_22_1/n53 ));
   CLKINVX1TS U2228 (.Y(\add_x_22_2/n121 ), 
	.A(\addr_calc/fir_read_calc/count[1] ));
   INVX2TS U2229 (.Y(n1972), 
	.A(\add_x_22_0/n84 ));
   CLKINVX1TS U2230 (.Y(\add_x_22_2/n105 ), 
	.A(FE_OFN245_addr_calc_fir_read_calc_count_5_));
   INVX1TS U2231 (.Y(\add_x_22_3/n19 ), 
	.A(\addr_calc/fir_write_calc/count[25] ));
   INVX2TS U2232 (.Y(n1970), 
	.A(\add_x_22_0/n80 ));
   INVX2TS U2234 (.Y(n1969), 
	.A(n1968));
   INVX2TS U2235 (.Y(n1840), 
	.A(n1839));
   CLKINVX2TS U2236 (.Y(n2553), 
	.A(\add_x_22_4/n105 ));
   INVX2TS U2237 (.Y(n1877), 
	.A(\add_x_22_3/n80 ));
   INVX2TS U2238 (.Y(n1974), 
	.A(n1973));
   CLKINVX1TS U2239 (.Y(\add_x_22_5/n114 ), 
	.A(\addr_calc/iir_write_calc/count[3] ));
   NOR2X1TS U2240 (.Y(\add_x_19_4/n48 ), 
	.B(FE_OFN351_offset_28_), 
	.A(\addr_calc/iir_read_calc/count[28] ));
   NOR2X4TS U2241 (.Y(\add_x_19_4/n97 ), 
	.B(FE_OFN384_offset_19_), 
	.A(\addr_calc/iir_read_calc/count[19] ));
   NOR2X4TS U2242 (.Y(\add_x_19_4/n58 ), 
	.B(\addr_calc/iir_read_calc/count[26] ), 
	.A(FE_OFN360_offset_26_));
   NOR2X1TS U2243 (.Y(\add_x_19_1/n78 ), 
	.B(FE_OCPUNCON1069_FE_OFN369_offset_23_), 
	.A(\addr_calc/fft_write_calc/count[23] ));
   NOR2X6TS U2244 (.Y(\add_x_19_1/n58 ), 
	.B(FE_OFN358_offset_26_), 
	.A(\addr_calc/fft_write_calc/count[26] ));
   NOR2X1TS U2245 (.Y(\add_x_19_1/n48 ), 
	.B(FE_OFN349_offset_28_), 
	.A(\addr_calc/fft_write_calc/count[28] ));
   NOR2X1TS U2246 (.Y(\add_x_19_1/n110 ), 
	.B(FE_OFN395_offset_16_), 
	.A(\addr_calc/fft_write_calc/count[16] ));
   NOR2X2TS U2247 (.Y(\add_x_19_2/n175 ), 
	.B(FE_OFN443_offset_4_), 
	.A(\addr_calc/fir_read_calc/count[4] ));
   NOR2X6TS U2248 (.Y(\add_x_19_5/n81 ), 
	.B(FE_OCPUNCON1877_FE_OFN374_offset_22_), 
	.A(\addr_calc/iir_write_calc/count[22] ));
   NOR2X4TS U2249 (.Y(\add_x_19_5/n58 ), 
	.B(FE_OFN360_offset_26_), 
	.A(\addr_calc/iir_write_calc/count[26] ));
   INVX2TS U2250 (.Y(n1679), 
	.A(\DP_OP_159_297_3515/n950 ));
   NOR2X2TS U2251 (.Y(\add_x_19_3/n58 ), 
	.B(FE_OFN359_offset_26_), 
	.A(FE_OFN267_addr_calc_fir_write_calc_count_26_));
   NOR2X2TS U2252 (.Y(\add_x_19_0/n48 ), 
	.B(FE_OFN352_offset_28_), 
	.A(\addr_calc/fft_read_calc/count[28] ));
   NOR2X2TS U2253 (.Y(\add_x_19_3/n66 ), 
	.B(FE_OFN368_offset_24_), 
	.A(\addr_calc/fir_write_calc/count[24] ));
   NOR2X1TS U2254 (.Y(\add_x_19_0/n58 ), 
	.B(FE_OFN359_offset_26_), 
	.A(\addr_calc/fft_read_calc/count[26] ));
   NOR2X4TS U2255 (.Y(\add_x_19_3/n78 ), 
	.B(FE_OFN371_offset_23_), 
	.A(\addr_calc/fir_write_calc/count[23] ));
   INVX2TS U2256 (.Y(n1680), 
	.A(n1641));
   INVX2TS U2257 (.Y(n1681), 
	.A(\DP_OP_159_297_3515/n873 ));
   OR2X1TS U2258 (.Y(n2630), 
	.B(FE_OFN339_offset_31_), 
	.A(FE_OFN262_addr_calc_fir_write_calc_count_31_));
   NOR2X1TS U2259 (.Y(\add_x_19_3/n110 ), 
	.B(FE_OFN396_offset_16_), 
	.A(\addr_calc/fir_write_calc/count[16] ));
   INVX2TS U2260 (.Y(n1682), 
	.A(\DP_OP_159_297_3515/n871 ));
   INVX2TS U2262 (.Y(\add_x_22_0/n89 ), 
	.A(\addr_calc/fft_read_calc/count[9] ));
   INVX2TS U2264 (.Y(n1850), 
	.A(\addr_calc/iir_write_calc/count[29] ));
   INVX2TS U2265 (.Y(\add_x_22_0/n92 ), 
	.A(\addr_calc/fft_read_calc/count[8] ));
   INVX2TS U2266 (.Y(\add_x_22_3/n30 ), 
	.A(\addr_calc/fir_write_calc/count[23] ));
   INVX2TS U2267 (.Y(n1973), 
	.A(\addr_calc/iir_write_calc/count[28] ));
   INVX2TS U2268 (.Y(\add_x_22_1/n74 ), 
	.A(\addr_calc/fft_write_calc/count[12] ));
   INVX2TS U2270 (.Y(n1685), 
	.A(n1907));
   INVX2TS U2272 (.Y(\add_x_22_0/n49 ), 
	.A(\addr_calc/fft_read_calc/count[18] ));
   INVX2TS U2273 (.Y(\add_x_22_4/n7 ), 
	.A(\addr_calc/iir_read_calc/count[28] ));
   INVX2TS U2274 (.Y(\add_x_22_1/n71 ), 
	.A(\addr_calc/fft_write_calc/count[13] ));
   INVX2TS U2275 (.Y(n1839), 
	.A(\addr_calc/iir_read_calc/count[29] ));
   INVX2TS U2276 (.Y(n1964), 
	.A(\addr_calc/iir_write_calc/count[23] ));
   INVX2TS U2277 (.Y(\add_x_22_0/n84 ), 
	.A(\addr_calc/fft_read_calc/count[10] ));
   INVX3TS U2278 (.Y(n1687), 
	.A(n1923));
   INVX2TS U2279 (.Y(\add_x_22_0/n80 ), 
	.A(\addr_calc/fft_read_calc/count[11] ));
   INVX2TS U2280 (.Y(\add_x_22_1/n53 ), 
	.A(\addr_calc/fft_write_calc/count[17] ));
   INVX2TS U2281 (.Y(n1957), 
	.A(\addr_calc/iir_write_calc/count[19] ));
   INVX2TS U2282 (.Y(n2050), 
	.A(\addr_calc/iir_write_calc/count[24] ));
   INVX2TS U2283 (.Y(n1919), 
	.A(\addr_calc/iir_read_calc/count[17] ));
   INVX2TS U2284 (.Y(\add_x_22_3/n80 ), 
	.A(\addr_calc/fir_write_calc/count[11] ));
   INVX2TS U2285 (.Y(\add_x_22_3/n105 ), 
	.A(\addr_calc/fir_write_calc/count[5] ));
   INVX2TS U2286 (.Y(n1688), 
	.A(n1971));
   INVX2TS U2287 (.Y(\add_x_22_4/n30 ), 
	.A(\addr_calc/iir_read_calc/count[23] ));
   INVX2TS U2289 (.Y(\add_x_22_4/n71 ), 
	.A(\addr_calc/iir_read_calc/count[13] ));
   INVX2TS U2290 (.Y(n2065), 
	.A(n2814));
   INVX2TS U2291 (.Y(n2062), 
	.A(n2815));
   INVX2TS U2292 (.Y(n2786), 
	.A(\addr_calc/iir_read_calc/count[0] ));
   INVX2TS U2293 (.Y(n2791), 
	.A(\addr_calc/iir_write_calc/count[0] ));
   INVX2TS U2294 (.Y(\add_x_22_4/n92 ), 
	.A(\addr_calc/iir_read_calc/count[8] ));
   INVX2TS U2295 (.Y(\add_x_22_1/n30 ), 
	.A(\addr_calc/fft_write_calc/count[23] ));
   INVX2TS U2296 (.Y(n2040), 
	.A(\addr_calc/fft_read_calc/count[22] ));
   INVX2TS U2297 (.Y(\add_x_22_1/n114 ), 
	.A(\addr_calc/fft_write_calc/count[3] ));
   INVX2TS U2298 (.Y(n1943), 
	.A(\addr_calc/fft_read_calc/count[27] ));
   INVX2TS U2299 (.Y(\add_x_22_0/n7 ), 
	.A(\addr_calc/fft_read_calc/count[28] ));
   INVX2TS U2300 (.Y(\add_x_22_1/n98 ), 
	.A(\addr_calc/fft_write_calc/count[7] ));
   INVX2TS U2302 (.Y(\add_x_22_1/n92 ), 
	.A(\addr_calc/fft_write_calc/count[8] ));
   INVX2TS U2303 (.Y(\add_x_22_1/n89 ), 
	.A(\addr_calc/fft_write_calc/count[9] ));
   INVX2TS U2304 (.Y(\add_x_22_1/n84 ), 
	.A(\addr_calc/fft_write_calc/count[10] ));
   INVX2TS U2305 (.Y(\add_x_22_1/n15 ), 
	.A(\addr_calc/fft_write_calc/count[26] ));
   INVX2TS U2306 (.Y(\add_x_22_2/n53 ), 
	.A(\addr_calc/fir_read_calc/count[17] ));
   INVX2TS U2307 (.Y(\add_x_22_2/n114 ), 
	.A(\addr_calc/fir_read_calc/count[3] ));
   INVX2TS U2308 (.Y(\add_x_22_2/n92 ), 
	.A(\addr_calc/fir_read_calc/count[8] ));
   INVX2TS U2310 (.Y(\add_x_22_2/n109 ), 
	.A(\addr_calc/fir_read_calc/count[4] ));
   INVX2TS U2311 (.Y(\add_x_22_5/n89 ), 
	.A(\addr_calc/iir_write_calc/count[9] ));
   INVX2TS U2312 (.Y(\add_x_22_5/n15 ), 
	.A(\addr_calc/iir_write_calc/count[26] ));
   INVX2TS U2313 (.Y(\add_x_22_5/n80 ), 
	.A(\addr_calc/iir_write_calc/count[11] ));
   INVX2TS U2314 (.Y(\add_x_22_2/n46 ), 
	.A(\addr_calc/fir_read_calc/count[19] ));
   INVX2TS U2315 (.Y(\add_x_22_2/n64 ), 
	.A(\addr_calc/fir_read_calc/count[15] ));
   INVX2TS U2316 (.Y(\add_x_22_5/n92 ), 
	.A(\addr_calc/iir_write_calc/count[8] ));
   INVX2TS U2317 (.Y(\add_x_22_2/n74 ), 
	.A(\addr_calc/fir_read_calc/count[12] ));
   INVX2TS U2318 (.Y(\add_x_22_2/n80 ), 
	.A(\addr_calc/fir_read_calc/count[11] ));
   INVX2TS U2319 (.Y(\add_x_22_3/n98 ), 
	.A(\addr_calc/fir_write_calc/count[7] ));
   INVX2TS U2321 (.Y(\add_x_22_3/n89 ), 
	.A(\addr_calc/fir_write_calc/count[9] ));
   INVX2TS U2322 (.Y(n1691), 
	.A(n1981));
   INVX2TS U2323 (.Y(\add_x_22_1/n7 ), 
	.A(\addr_calc/fft_write_calc/count[28] ));
   INVX2TS U2324 (.Y(\add_x_22_5/n57 ), 
	.A(\addr_calc/iir_write_calc/count[16] ));
   INVX2TS U2325 (.Y(n1930), 
	.A(\addr_calc/fft_write_calc/count[11] ));
   INVX2TS U2326 (.Y(n1852), 
	.A(\addr_calc/fft_write_calc/count[29] ));
   INVX2TS U2327 (.Y(n1982), 
	.A(\addr_calc/fir_read_calc/count[24] ));
   INVX2TS U2329 (.Y(\add_x_22_5/n84 ), 
	.A(\addr_calc/iir_write_calc/count[10] ));
   INVX2TS U2330 (.Y(n1834), 
	.A(\addr_calc/fir_write_calc/count[27] ));
   INVX2TS U2331 (.Y(\add_x_22_5/n121 ), 
	.A(\addr_calc/iir_write_calc/count[1] ));
   INVX2TS U2332 (.Y(\add_x_22_3/n7 ), 
	.A(\addr_calc/fir_write_calc/count[28] ));
   INVX2TS U2333 (.Y(\add_x_22_3/n71 ), 
	.A(\addr_calc/fir_write_calc/count[13] ));
   INVX2TS U2334 (.Y(\add_x_22_2/n71 ), 
	.A(\addr_calc/fir_read_calc/count[13] ));
   CLKINVX2TS U2338 (.Y(n2504), 
	.A(n2503));
   CLKINVX2TS U2339 (.Y(n2502), 
	.A(n2501));
   CLKINVX2TS U2340 (.Y(n2506), 
	.A(n2505));
   CLKINVX2TS U2344 (.Y(n2352), 
	.A(n2351));
   CLKINVX2TS U2349 (.Y(n2356), 
	.A(n2355));
   CLKINVX2TS U2352 (.Y(n2518), 
	.A(n2517));
   CLKINVX2TS U2354 (.Y(n2520), 
	.A(n2519));
   CLKINVX2TS U2356 (.Y(n2534), 
	.A(n2533));
   CLKINVX2TS U2362 (.Y(n2536), 
	.A(n2535));
   CLKINVX2TS U2366 (.Y(n2540), 
	.A(n2539));
   CLKINVX2TS U2372 (.Y(n2346), 
	.A(n2345));
   CLKINVX2TS U2375 (.Y(n2510), 
	.A(n2509));
   CLKINVX2TS U2377 (.Y(n2526), 
	.A(n2525));
   CLKINVX2TS U2381 (.Y(n2542), 
	.A(n2541));
   CLKINVX2TS U2384 (.Y(n2548), 
	.A(n2547));
   CLKINVX2TS U2385 (.Y(n2350), 
	.A(n2349));
   CLKINVX2TS U2387 (.Y(n2532), 
	.A(n2531));
   CLKINVX2TS U2389 (.Y(n2516), 
	.A(n2515));
   CLKINVX2TS U2392 (.Y(n2358), 
	.A(n2357));
   CLKINVX2TS U2393 (.Y(n2512), 
	.A(n2511));
   CLKINVX2TS U2395 (.Y(n2546), 
	.A(n2545));
   CLKINVX2TS U2398 (.Y(n2530), 
	.A(n2529));
   CLKINVX2TS U2399 (.Y(n2528), 
	.A(n2527));
   CLKINVX2TS U2401 (.Y(n2514), 
	.A(n2513));
   CLKINVX2TS U2402 (.Y(n2354), 
	.A(n2353));
   CLKINVX2TS U2405 (.Y(n2522), 
	.A(n2521));
   CLKINVX2TS U2407 (.Y(n2538), 
	.A(n2537));
   CLKINVX2TS U2410 (.Y(n2348), 
	.A(n2347));
   CLKINVX2TS U2412 (.Y(n2508), 
	.A(n2507));
   CLKINVX2TS U2416 (.Y(n2524), 
	.A(n2523));
   CLKINVX2TS U2420 (.Y(n2544), 
	.A(n2543));
   INVX2TS U2507 (.Y(n2325), 
	.A(n2324));
   CLKINVX2TS U2518 (.Y(n2360), 
	.A(n2359));
   XOR2X1TS U2547 (.Y(n2615), 
	.B(FE_OFN481_filesize_16_), 
	.A(\DP_OP_159_297_3515/n989 ));
   AO22X1TS U2548 (.Y(n1116), 
	.B1(\addr_calc/fir_write_calc/count[14] ), 
	.B0(FE_OCPUNCON1084_n2805), 
	.A1(\addr_calc/fir_write_calc/counter/N57 ), 
	.A0(FE_OFN48_n2803));
   INVX2TS U2549 (.Y(n1947), 
	.A(n1946));
   NOR2X2TS U2550 (.Y(\DP_OP_158_296_6262/n320 ), 
	.B(\DP_OP_158_296_6262/n329 ), 
	.A(\DP_OP_158_296_6262/n322 ));
   NOR2BX1TS U2553 (.Y(\DP_OP_159_297_3515/n648 ), 
	.B(\DP_OP_159_297_3515/n650 ), 
	.AN(n1692));
   XOR2X1TS U2554 (.Y(n1692), 
	.B(FE_OFN230_addr_calc_iir_write_calc_count_15_), 
	.A(n2616));
   OAI21X2TS U2555 (.Y(\add_x_19_4/n57 ), 
	.B0(\add_x_19_4/n59 ), 
	.A1(\add_x_19_4/n58 ), 
	.A0(\add_x_19_4/n60 ));
   AOI21X4TS U2556 (.Y(\add_x_19_4/n60 ), 
	.B0(\add_x_19_4/n62 ), 
	.A1(\add_x_19_4/n61 ), 
	.A0(\add_x_19_4/n69 ));
   NOR2X1TS U2557 (.Y(\DP_OP_159_297_3515/n623 ), 
	.B(\DP_OP_159_297_3515/n638 ), 
	.A(\DP_OP_159_297_3515/n625 ));
   NOR2X2TS U2558 (.Y(\DP_OP_159_297_3515/n587 ), 
	.B(\DP_OP_159_297_3515/n646 ), 
	.A(\DP_OP_159_297_3515/n589 ));
   NAND2X2TS U2559 (.Y(\DP_OP_159_297_3515/n589 ), 
	.B(\DP_OP_159_297_3515/n623 ), 
	.A(\DP_OP_159_297_3515/n591 ));
   XNOR2X1TS U2560 (.Y(\DP_OP_159_297_3515/n730 ), 
	.B(n2041), 
	.A(n2622));
   AO22X1TS U2561 (.Y(n1108), 
	.B1(\addr_calc/fir_write_calc/count[22] ), 
	.B0(FE_OCPUNCON1087_n2805), 
	.A1(\addr_calc/fir_write_calc/counter/N65 ), 
	.A0(n1762));
   NOR2X2TS U2562 (.Y(\add_x_19_3/n63 ), 
	.B(FE_OFN363_offset_25_), 
	.A(FE_OFN231_addr_calc_fir_write_calc_count_25_));
   NOR2X2TS U2563 (.Y(\DP_OP_158_296_6262/n131 ), 
	.B(\DP_OP_158_296_6262/n133 ), 
	.A(\DP_OP_158_296_6262/n148 ));
   NOR2X4TS U2565 (.Y(\DP_OP_159_297_3515/n688 ), 
	.B(\DP_OP_159_297_3515/n690 ), 
	.A(FE_OFN535_DP_OP_159_297_3515_n726));
   AND2X4TS U2566 (.Y(n1780), 
	.B(\DP_OP_159_297_3515/n688 ), 
	.A(\DP_OP_159_297_3515/n587 ));
   NAND2X2TS U2567 (.Y(\DP_OP_159_297_3515/n913 ), 
	.B(\DP_OP_159_297_3515/n914 ), 
	.A(FE_OCPUNCON1565_n1789));
   NOR2X1TS U2568 (.Y(\DP_OP_158_296_6262/n1855 ), 
	.B(n1664), 
	.A(\DP_OP_158_296_6262/n1863 ));
   AO22X4TS U2569 (.Y(n1128), 
	.B1(n1990), 
	.B0(FE_OCPUNCON1093_n2805), 
	.A1(\addr_calc/fir_write_calc/counter/N45 ), 
	.A0(FE_OFN51_n2803));
   NAND2X1TS U2571 (.Y(\DP_OP_159_297_3515/n934 ), 
	.B(\DP_OP_159_297_3515/n935 ), 
	.A(n1792));
   XNOR2X4TS U2572 (.Y(\addr_calc/iir_read_addr[19] ), 
	.B(\add_x_19_4/n13 ), 
	.A(\add_x_19_4/n99 ));
   INVX2TS U2573 (.Y(\add_x_22_5/n71 ), 
	.A(\addr_calc/iir_write_calc/count[13] ));
   XOR2X4TS U2574 (.Y(n1697), 
	.B(\DP_OP_158_296_6262/n1897 ), 
	.A(n1698));
   NOR4XLTS U2575 (.Y(n906), 
	.D(n908), 
	.C(n907), 
	.B(instruction[11]), 
	.A(instruction[12]));
   XOR2X4TS U2576 (.Y(n1699), 
	.B(n1679), 
	.A(\DP_OP_159_297_3515/n955 ));
   AO22X1TS U2577 (.Y(n1089), 
	.B1(\addr_calc/fir_read_calc/count[9] ), 
	.B0(FE_OFN63_n2809), 
	.A1(\addr_calc/fir_read_calc/counter/N52 ), 
	.A0(FE_OFN54_n2807));
   AO22X1TS U2578 (.Y(n1078), 
	.B1(\addr_calc/fir_read_calc/count[20] ), 
	.B0(FE_OFN66_n2809), 
	.A1(\addr_calc/fir_read_calc/counter/N63 ), 
	.A0(FE_OFN56_n2807));
   NOR2X1TS U2579 (.Y(\DP_OP_159_297_3515/n672 ), 
	.B(\DP_OP_159_297_3515/n674 ), 
	.A(\DP_OP_159_297_3515/n685 ));
   AO22X1TS U2580 (.Y(n1006), 
	.B1(n2559), 
	.B0(FE_OFN13_n2794), 
	.A1(\addr_calc/fft_read_calc/counter/N71 ), 
	.A0(FE_OFN4_n1755));
   AO22X2TS U2581 (.Y(n1027), 
	.B1(n1666), 
	.B0(FE_OFN16_n2794), 
	.A1(\addr_calc/fft_read_calc/counter/N50 ), 
	.A0(FE_OFN550_n1750));
   XNOR2X1TS U2582 (.Y(\DP_OP_159_297_3515/n685 ), 
	.B(n1945), 
	.A(n2618));
   AO22X1TS U2583 (.Y(n1014), 
	.B1(n2572), 
	.B0(FE_OFN11_n2794), 
	.A1(\addr_calc/fft_read_calc/counter/N63 ), 
	.A0(FE_OFN551_n1751));
   INVX2TS U2584 (.Y(n1792), 
	.A(n1782));
   AO22X1TS U2585 (.Y(n1021), 
	.B1(\addr_calc/fft_read_calc/count[13] ), 
	.B0(FE_OFN8_n2794), 
	.A1(\addr_calc/fft_read_calc/counter/N56 ), 
	.A0(FE_OFN6_n1750));
   AO22X1TS U2586 (.Y(n1020), 
	.B1(\addr_calc/fft_read_calc/count[14] ), 
	.B0(FE_OFN7_n2794), 
	.A1(\addr_calc/fft_read_calc/counter/N57 ), 
	.A0(n1755));
   AO22X1TS U2588 (.Y(n1022), 
	.B1(\addr_calc/fft_read_calc/count[12] ), 
	.B0(FE_OFN8_n2794), 
	.A1(\addr_calc/fft_read_calc/counter/N55 ), 
	.A0(FE_OFN1_n1751));
   AO22X1TS U2589 (.Y(n1012), 
	.B1(\addr_calc/fft_read_calc/count[22] ), 
	.B0(FE_OFN11_n2794), 
	.A1(\addr_calc/fft_read_calc/counter/N65 ), 
	.A0(FE_OFN552_n1751));
   XNOR2X4TS U2590 (.Y(n1702), 
	.B(n1678), 
	.A(\DP_OP_159_297_3515/n913 ));
   AO22X1TS U2591 (.Y(n1112), 
	.B1(\addr_calc/fir_write_calc/count[18] ), 
	.B0(FE_OCPUNCON1086_n2805), 
	.A1(\addr_calc/fir_write_calc/counter/N61 ), 
	.A0(FE_OFN49_n2803));
   XNOR2X4TS U2593 (.Y(n1703), 
	.B(\DP_OP_159_297_3515/n862 ), 
	.A(\DP_OP_159_297_3515/n948 ));
   AND2X8TS U2594 (.Y(n1715), 
	.B(\DP_OP_158_296_6262/n3 ), 
	.A(\DP_OP_158_296_6262/n62 ));
   XNOR2X1TS U2596 (.Y(\DP_OP_158_296_6262/n133 ), 
	.B(n2558), 
	.A(n1731));
   NOR2X1TS U2598 (.Y(\DP_OP_159_297_3515/n712 ), 
	.B(\DP_OP_159_297_3515/n723 ), 
	.A(\DP_OP_159_297_3515/n714 ));
   NAND2X8TS U2609 (.Y(\addr_calc/fir_read_calc/counter/N38 ), 
	.B(n1716), 
	.A(n1715));
   AND2X4TS U2610 (.Y(n1716), 
	.B(\DP_OP_158_296_6262/n280 ), 
	.A(\DP_OP_158_296_6262/n179 ));
   NAND2X2TS U2611 (.Y(\DP_OP_159_297_3515/n906 ), 
	.B(FE_OCPUNCON1566_n1789), 
	.A(\DP_OP_159_297_3515/n907 ));
   XOR2X1TS U2612 (.Y(n2618), 
	.B(n1682), 
	.A(\DP_OP_159_297_3515/n1010 ));
   NOR2X2TS U2613 (.Y(\DP_OP_158_296_6262/n1833 ), 
	.B(\DP_OP_158_296_6262/n1834 ), 
	.A(FE_OCPUNCON1567_n1717));
   NAND2X1TS U2614 (.Y(\DP_OP_159_297_3515/n996 ), 
	.B(\DP_OP_159_297_3515/n997 ), 
	.A(n1788));
   OR2X2TS U2615 (.Y(n1728), 
	.B(\DP_OP_158_296_6262/n1987 ), 
	.A(\DP_OP_158_296_6262/n2011 ));
   AO22X1TS U2616 (.Y(n1111), 
	.B1(n1670), 
	.B0(FE_OCPUNCON1086_n2805), 
	.A1(\addr_calc/fir_write_calc/counter/N62 ), 
	.A0(n1762));
   AO22X1TS U2617 (.Y(n1056), 
	.B1(n1932), 
	.B0(FE_OCPN1911_FE_OFN17_n2797), 
	.A1(\addr_calc/fft_write_calc/counter/N53 ), 
	.A0(n2795));
   AO22X1TS U2618 (.Y(n1057), 
	.B1(n1934), 
	.B0(FE_OFN19_n2797), 
	.A1(\addr_calc/fft_write_calc/counter/N52 ), 
	.A0(FE_OFN28_n2795));
   AO22X4TS U2619 (.Y(n1059), 
	.B1(n1936), 
	.B0(FE_OFN26_n2797), 
	.A1(\addr_calc/fft_write_calc/counter/N50 ), 
	.A0(FE_OFN35_n2795));
   AO22X1TS U2620 (.Y(n1051), 
	.B1(n1976), 
	.B0(FE_OFN18_n2797), 
	.A1(\addr_calc/fft_write_calc/counter/N58 ), 
	.A0(FE_OFN27_n2795));
   XNOR2X4TS U2621 (.Y(n1731), 
	.B(FE_OFN473_filesize_23_), 
	.A(\DP_OP_158_296_6262/n1881 ));
   AO22X1TS U2623 (.Y(n1045), 
	.B1(\addr_calc/fft_write_calc/count[21] ), 
	.B0(FE_OFN21_n2797), 
	.A1(\addr_calc/fft_write_calc/counter/N64 ), 
	.A0(FE_OFN30_n2795));
   AO22X1TS U2624 (.Y(n1047), 
	.B1(\addr_calc/fft_write_calc/count[19] ), 
	.B0(FE_OFN20_n2797), 
	.A1(\addr_calc/fft_write_calc/counter/N62 ), 
	.A0(FE_OFN29_n2795));
   XNOR2X1TS U2625 (.Y(n2616), 
	.B(\DP_OP_159_297_3515/n869 ), 
	.A(\DP_OP_159_297_3515/n996 ));
   NAND2X1TS U2626 (.Y(\DP_OP_159_297_3515/n1003 ), 
	.B(\DP_OP_159_297_3515/n1004 ), 
	.A(n1787));
   AO22X1TS U2630 (.Y(n1053), 
	.B1(n1927), 
	.B0(FE_OFN18_n2797), 
	.A1(\addr_calc/fft_write_calc/counter/N56 ), 
	.A0(FE_OFN27_n2795));
   AO22X1TS U2631 (.Y(n1054), 
	.B1(n2023), 
	.B0(FE_OCPN1911_FE_OFN17_n2797), 
	.A1(\addr_calc/fft_write_calc/counter/N55 ), 
	.A0(n2795));
   AO22X1TS U2634 (.Y(n1076), 
	.B1(\addr_calc/fir_read_calc/count[22] ), 
	.B0(FE_OFN67_n2809), 
	.A1(\addr_calc/fir_read_calc/counter/N65 ), 
	.A0(FE_OFN57_n2807));
   CLKXOR2X8TS U2635 (.Y(n1775), 
	.B(n2330), 
	.A(\DP_OP_158_296_6262/n1847 ));
   MXI2X1TS U2636 (.Y(n1130), 
	.S0(n2805), 
	.B(\addr_calc/fir_write_calc/counter/N43 ), 
	.A(n2806));
   NOR2X4TS U2637 (.Y(n2787), 
	.B(n1737), 
	.A(n1781));
   XNOR2X1TS U2638 (.Y(\DP_OP_159_297_3515/n593 ), 
	.B(n2048), 
	.A(n1697));
   NAND2X1TS U2639 (.Y(\DP_OP_159_297_3515/n1017 ), 
	.B(\DP_OP_159_297_3515/n1018 ), 
	.A(n1787));
   NOR2X2TS U2640 (.Y(\DP_OP_159_297_3515/n591 ), 
	.B(\DP_OP_159_297_3515/n593 ), 
	.A(\DP_OP_159_297_3515/n610 ));
   NOR2X1TS U2641 (.Y(\DP_OP_158_296_6262/n102 ), 
	.B(\DP_OP_158_296_6262/n119 ), 
	.A(\DP_OP_158_296_6262/n104 ));
   NAND2X1TS U2643 (.Y(\DP_OP_159_297_3515/n989 ), 
	.B(\DP_OP_159_297_3515/n990 ), 
	.A(n1788));
   NOR2X1TS U2644 (.Y(\DP_OP_158_296_6262/n240 ), 
	.B(\DP_OP_158_296_6262/n242 ), 
	.A(\DP_OP_158_296_6262/n255 ));
   AO22X1TS U2646 (.Y(n952), 
	.B1(n2556), 
	.B0(FE_OFN91_n1192), 
	.A1(\addr_calc/iir_read_calc/counter/N62 ), 
	.A0(FE_OFN78_n2787));
   NOR2X2TS U2647 (.Y(\add_x_19_4/n131 ), 
	.B(FE_OCPUNCON1073_FE_OFN410_offset_12_), 
	.A(\addr_calc/iir_read_calc/count[12] ));
   AO22X1TS U2651 (.Y(n994), 
	.B1(n2041), 
	.B0(FE_OCPUNCON1568_n2812), 
	.A1(\addr_calc/iir_write_calc/counter/N51 ), 
	.A0(n2813));
   AO22X1TS U2652 (.Y(n960), 
	.B1(\addr_calc/iir_read_calc/count[11] ), 
	.B0(FE_OFN85_n2654), 
	.A1(\addr_calc/iir_read_calc/counter/N54 ), 
	.A0(n2787));
   AO22X1TS U2653 (.Y(n993), 
	.B1(n2562), 
	.B0(FE_OCPUNCON1568_n2812), 
	.A1(\addr_calc/iir_write_calc/counter/N52 ), 
	.A0(n2813));
   AO22X1TS U2656 (.Y(n951), 
	.B1(\addr_calc/iir_read_calc/count[20] ), 
	.B0(FE_OFN91_n1192), 
	.A1(\addr_calc/iir_read_calc/counter/N63 ), 
	.A0(FE_OFN79_n2787));
   AO22X1TS U2657 (.Y(n1075), 
	.B1(n2558), 
	.B0(FE_OFN67_n2809), 
	.A1(\addr_calc/fir_read_calc/counter/N66 ), 
	.A0(FE_OFN57_n2807));
   NOR2X2TS U2659 (.Y(\DP_OP_158_296_6262/n1826 ), 
	.B(\DP_OP_158_296_6262/n1827 ), 
	.A(FE_OCPUNCON1567_n1717));
   XNOR2X4TS U2660 (.Y(n1756), 
	.B(n2368), 
	.A(\DP_OP_158_296_6262/n1957 ));
   NOR2X1TS U2661 (.Y(\DP_OP_158_296_6262/n1957 ), 
	.B(n1455), 
	.A(n1693));
   INVX2TS U2662 (.Y(n1785), 
	.A(\add_x_22_4/n74 ));
   NAND2X2TS U2663 (.Y(\add_x_19_4/n132 ), 
	.B(FE_OCPUNCON1073_FE_OFN410_offset_12_), 
	.A(\addr_calc/iir_read_calc/count[12] ));
   XNOR2X1TS U2664 (.Y(\DP_OP_158_296_6262/n87 ), 
	.B(FE_OFN270_addr_calc_fir_read_calc_count_26_), 
	.A(\DP_OP_158_296_6262/n833 ));
   NOR2X2TS U2665 (.Y(\DP_OP_158_296_6262/n179 ), 
	.B(\DP_OP_158_296_6262/n238 ), 
	.A(\DP_OP_158_296_6262/n181 ));
   NAND2X1TS U2666 (.Y(\DP_OP_158_296_6262/n238 ), 
	.B(\DP_OP_158_296_6262/n240 ), 
	.A(\DP_OP_158_296_6262/n264 ));
   NAND2X2TS U2667 (.Y(\DP_OP_158_296_6262/n181 ), 
	.B(\DP_OP_158_296_6262/n215 ), 
	.A(\DP_OP_158_296_6262/n183 ));
   NOR2X1TS U2668 (.Y(\DP_OP_158_296_6262/n183 ), 
	.B(\DP_OP_158_296_6262/n185 ), 
	.A(\DP_OP_158_296_6262/n202 ));
   INVX2TS U2670 (.Y(\DP_OP_158_296_6262/n838 ), 
	.A(\DP_OP_158_296_6262/n2051 ));
   XNOR2X1TS U2671 (.Y(\DP_OP_158_296_6262/n217 ), 
	.B(n1884), 
	.A(n1729));
   AO22X1TS U2672 (.Y(n1058), 
	.B1(n2026), 
	.B0(FE_OFN19_n2797), 
	.A1(\addr_calc/fft_write_calc/counter/N51 ), 
	.A0(FE_OFN28_n2795));
   AO22X1TS U2673 (.Y(n1043), 
	.B1(n2555), 
	.B0(FE_OFN21_n2797), 
	.A1(\addr_calc/fft_write_calc/counter/N66 ), 
	.A0(FE_OFN30_n2795));
   AO22X1TS U2674 (.Y(n1038), 
	.B1(n2557), 
	.B0(FE_OFN22_n2797), 
	.A1(\addr_calc/fft_write_calc/counter/N71 ), 
	.A0(FE_OFN31_n2795));
   AO22X4TS U2676 (.Y(n1063), 
	.B1(n2568), 
	.B0(FE_OFN25_n2797), 
	.A1(\addr_calc/fft_write_calc/counter/N46 ), 
	.A0(FE_OFN34_n2795));
   XNOR2X1TS U2679 (.Y(\DP_OP_159_297_3515/n694 ), 
	.B(n2044), 
	.A(n2619));
   XNOR2X4TS U2680 (.Y(n2619), 
	.B(\DP_OP_158_296_6262/n1952 ), 
	.A(\DP_OP_159_297_3515/n1017 ));
   NAND2X2TS U2681 (.Y(\DP_OP_158_296_6262/n18 ), 
	.B(n1653), 
	.A(\DP_OP_158_296_6262/n37 ));
   XNOR2X1TS U2682 (.Y(\DP_OP_158_296_6262/n104 ), 
	.B(\addr_calc/fir_read_calc/count[25] ), 
	.A(n1655));
   XNOR2X1TS U2683 (.Y(\DP_OP_158_296_6262/n119 ), 
	.B(n1983), 
	.A(FE_OCPN1732_n1718));
   AND4X1TS U2684 (.Y(n817), 
	.D(\add_x_22_4/n71 ), 
	.C(\add_x_22_4/n67 ), 
	.B(\add_x_22_4/n64 ), 
	.A(\add_x_22_4/n57 ));
   INVX2TS U2685 (.Y(\add_x_22_4/n64 ), 
	.A(\addr_calc/iir_read_calc/count[15] ));
   NAND2X2TS U2686 (.Y(\DP_OP_159_297_3515/n920 ), 
	.B(FE_OCPUNCON1565_n1789), 
	.A(\DP_OP_159_297_3515/n921 ));
   XNOR2X1TS U2687 (.Y(\DP_OP_158_296_6262/n185 ), 
	.B(n1881), 
	.A(n1654));
   CLKXOR2X4TS U2688 (.Y(n2595), 
	.B(FE_OFN495_filesize_5_), 
	.A(\DP_OP_158_296_6262/n2004 ));
   XNOR2X4TS U2689 (.Y(\addr_calc/iir_read_addr[27] ), 
	.B(\add_x_19_4/n5 ), 
	.A(\add_x_19_4/n57 ));
   XOR2X4TS U2690 (.Y(\DP_OP_158_296_6262/n2060 ), 
	.B(n2341), 
	.A(\DP_OP_158_296_6262/n1833 ));
   NOR2X1TS U2691 (.Y(\DP_OP_158_296_6262/n215 ), 
	.B(\DP_OP_158_296_6262/n230 ), 
	.A(\DP_OP_158_296_6262/n217 ));
   AO22X1TS U2692 (.Y(n959), 
	.B1(n1785), 
	.B0(n1192), 
	.A1(\addr_calc/iir_read_calc/counter/N55 ), 
	.A0(FE_OCPUNCON1878_n2787));
   AO22X1TS U2693 (.Y(n957), 
	.B1(n1784), 
	.B0(n1192), 
	.A1(\addr_calc/iir_read_calc/counter/N57 ), 
	.A0(FE_OCPUNCON1880_n2787));
   NOR2X2TS U2694 (.Y(\DP_OP_158_296_6262/n1991 ), 
	.B(n2366), 
	.A(\DP_OP_158_296_6262/n1998 ));
   NAND2X1TS U2695 (.Y(\DP_OP_159_297_3515/n852 ), 
	.B(\DP_OP_159_297_3515/n930 ), 
	.A(\DP_OP_159_297_3515/n956 ));
   NOR2X1TS U2696 (.Y(\DP_OP_158_296_6262/n1916 ), 
	.B(\DP_OP_158_296_6262/n1917 ), 
	.A(n2589));
   NAND2X2TS U2697 (.Y(\DP_OP_158_296_6262/n64 ), 
	.B(\DP_OP_158_296_6262/n102 ), 
	.A(\DP_OP_158_296_6262/n66 ));
   NAND2X2TS U2698 (.Y(\DP_OP_158_296_6262/n129 ), 
	.B(\DP_OP_158_296_6262/n131 ), 
	.A(\DP_OP_158_296_6262/n159 ));
   NOR2X1TS U2700 (.Y(\DP_OP_158_296_6262/n1909 ), 
	.B(\DP_OP_158_296_6262/n1910 ), 
	.A(n2589));
   NOR2X1TS U2701 (.Y(\DP_OP_158_296_6262/n1943 ), 
	.B(\DP_OP_158_296_6262/n1944 ), 
	.A(n1728));
   XOR2X1TS U2702 (.Y(\DP_OP_158_296_6262/n2051 ), 
	.B(n1679), 
	.A(\DP_OP_158_296_6262/n1895 ));
   AOI21X4TS U2703 (.Y(n2809), 
	.B0(FE_OFN562_n2060), 
	.A1(FE_OFN330_data_to_fir), 
	.A0(\addr_calc/fir_read_calc/counter/N38 ));
   XOR2X4TS U2704 (.Y(\DP_OP_158_296_6262/n2048 ), 
	.B(FE_OFN479_filesize_18_), 
	.A(\DP_OP_158_296_6262/n1916 ));
   NAND2X1TS U2707 (.Y(\DP_OP_159_297_3515/n690 ), 
	.B(\DP_OP_159_297_3515/n712 ), 
	.A(\DP_OP_159_297_3515/n692 ));
   NOR2X1TS U2708 (.Y(\DP_OP_159_297_3515/n692 ), 
	.B(\DP_OP_159_297_3515/n694 ), 
	.A(\DP_OP_159_297_3515/n705 ));
   XNOR2X4TS U2709 (.Y(n2621), 
	.B(\DP_OP_158_296_6262/n1966 ), 
	.A(\DP_OP_159_297_3515/n1031 ));
   AO22X1TS U2710 (.Y(n980), 
	.B1(n2579), 
	.B0(FE_OCPUNCON1572_n2812), 
	.A1(\addr_calc/iir_write_calc/counter/N65 ), 
	.A0(FE_OCPUNCON1883_n2813));
   AO22X1TS U2711 (.Y(n1070), 
	.B1(\addr_calc/fir_read_calc/count[28] ), 
	.B0(FE_OFN67_n2809), 
	.A1(\addr_calc/fir_read_calc/counter/N71 ), 
	.A0(FE_OFN57_n2807));
   MXI2X1TS U2712 (.Y(n1002), 
	.S0(FE_OCPUNCON1569_n2812), 
	.B(n2791), 
	.A(n2792));
   XOR2X4TS U2713 (.Y(\DP_OP_159_297_3515/n1128 ), 
	.B(\DP_OP_158_296_6262/n1911 ), 
	.A(\DP_OP_159_297_3515/n976 ));
   MXI2X1TS U2715 (.Y(n1098), 
	.S0(FE_OFN64_n2809), 
	.B(n2810), 
	.A(n2811));
   AO22X1TS U2716 (.Y(n1004), 
	.B1(\addr_calc/fft_read_calc/count[30] ), 
	.B0(FE_OFN14_n2794), 
	.A1(\addr_calc/fft_read_calc/counter/N73 ), 
	.A0(FE_OFN551_n1751));
   NAND2X1TS U2731 (.Y(\DP_OP_159_297_3515/n971 ), 
	.B(FE_OFN479_filesize_18_), 
	.A(FE_OFN480_filesize_17_));
   INVXLTS U2732 (.Y(\DP_OP_159_297_3515/n964 ), 
	.A(FE_OFN478_filesize_19_));
   AO22X1TS U2734 (.Y(n1036), 
	.B1(\addr_calc/fft_write_calc/count[30] ), 
	.B0(FE_OFN24_n2797), 
	.A1(\addr_calc/fft_write_calc/counter/N73 ), 
	.A0(FE_OFN33_n2795));
   AO22X1TS U2735 (.Y(n1069), 
	.B1(\addr_calc/fir_read_calc/count[29] ), 
	.B0(FE_OFN69_n2809), 
	.A1(\addr_calc/fir_read_calc/counter/N72 ), 
	.A0(FE_OFN59_n2807));
   INVX2TS U2736 (.Y(\DP_OP_159_297_3515/n957 ), 
	.A(\DP_OP_159_297_3515/n956 ));
   AO22X1TS U2737 (.Y(n1084), 
	.B1(\addr_calc/fir_read_calc/count[14] ), 
	.B0(n2809), 
	.A1(\addr_calc/fir_read_calc/counter/N57 ), 
	.A0(FE_OFN52_n2807));
   NOR2X1TS U2739 (.Y(\DP_OP_159_297_3515/n930 ), 
	.B(\DP_OP_159_297_3515/n931 ), 
	.A(\DP_OP_159_297_3515/n943 ));
   AO22X1TS U2740 (.Y(n953), 
	.B1(\addr_calc/iir_read_calc/count[18] ), 
	.B0(FE_OFN90_n1192), 
	.A1(\addr_calc/iir_read_calc/counter/N61 ), 
	.A0(FE_OFN78_n2787));
   NOR2X2TS U2741 (.Y(\add_x_19_0/n165 ), 
	.B(FE_OCPUNCON726_FE_OFN435_offset_6_), 
	.A(FE_OFN225_addr_calc_fft_read_calc_count_6_));
   NOR2X6TS U2742 (.Y(\add_x_19_4/n78 ), 
	.B(\addr_calc/iir_read_calc/count[23] ), 
	.A(FE_OFN372_offset_23_));
   INVX2TS U2751 (.Y(n1860), 
	.A(n2815));
   INVX2TS U2752 (.Y(\add_x_22_3/n114 ), 
	.A(\addr_calc/fir_write_calc/count[3] ));
   NOR2X1TS U2754 (.Y(\add_x_19_2/n55 ), 
	.B(FE_OFN354_offset_27_), 
	.A(\addr_calc/fir_read_calc/count[27] ));
   INVX2TS U2755 (.Y(\add_x_22_3/n84 ), 
	.A(\addr_calc/fir_write_calc/count[10] ));
   INVX2TS U2756 (.Y(n1875), 
	.A(\addr_calc/fir_read_calc/count[25] ));
   INVX2TS U2757 (.Y(n1876), 
	.A(n1875));
   INVX2TS U2758 (.Y(n1882), 
	.A(\addr_calc/fir_write_calc/count[15] ));
   INVX2TS U2759 (.Y(n1885), 
	.A(\addr_calc/fir_write_calc/count[17] ));
   INVX2TS U2760 (.Y(n1886), 
	.A(n1885));
   INVX2TS U2761 (.Y(n1887), 
	.A(\addr_calc/fir_read_calc/count[16] ));
   NOR4XLTS U2762 (.Y(n864), 
	.D(\addr_calc/fir_write_calc/count[28] ), 
	.C(FE_OFN273_addr_calc_fir_write_calc_count_29_), 
	.B(\addr_calc/fir_write_calc/count[2] ), 
	.A(FE_OFN238_addr_calc_fir_write_calc_count_30_));
   INVX2TS U2763 (.Y(n1898), 
	.A(\add_x_22_4/n121 ));
   INVX2TS U2764 (.Y(\add_x_22_4/n121 ), 
	.A(\addr_calc/iir_read_calc/count[1] ));
   INVX2TS U2766 (.Y(n1912), 
	.A(\addr_calc/fft_write_calc/count[27] ));
   INVX2TS U2767 (.Y(n1913), 
	.A(n1912));
   INVX2TS U2768 (.Y(n1914), 
	.A(\addr_calc/fft_write_calc/count[25] ));
   INVX2TS U2769 (.Y(n1915), 
	.A(n1914));
   INVX2TS U2770 (.Y(n1917), 
	.A(\addr_calc/fft_write_calc/count[21] ));
   INVX2TS U2771 (.Y(n1922), 
	.A(n1921));
   INVX2TS U2772 (.Y(n1926), 
	.A(n1925));
   INVX2TS U2774 (.Y(n1931), 
	.A(\add_x_22_5/n121 ));
   INVX2TS U2775 (.Y(\add_x_22_5/n109 ), 
	.A(\addr_calc/iir_write_calc/count[4] ));
   INVX2TS U2776 (.Y(n1939), 
	.A(\add_x_22_1/n109 ));
   AO22X4TS U2777 (.Y(n1062), 
	.B1(n1939), 
	.B0(FE_OFN26_n2797), 
	.A1(\addr_calc/fft_write_calc/counter/N47 ), 
	.A0(FE_OFN35_n2795));
   INVX2TS U2778 (.Y(\add_x_22_1/n109 ), 
	.A(\addr_calc/fft_write_calc/count[4] ));
   INVX2TS U2779 (.Y(n1941), 
	.A(\add_x_22_1/n121 ));
   INVX2TS U2780 (.Y(\add_x_22_1/n121 ), 
	.A(\addr_calc/fft_write_calc/count[1] ));
   INVX2TS U2781 (.Y(n1946), 
	.A(\addr_calc/fft_read_calc/count[25] ));
   INVX2TS U2782 (.Y(n1949), 
	.A(\addr_calc/fft_read_calc/count[23] ));
   INVX2TS U2783 (.Y(n1950), 
	.A(n1949));
   INVX2TS U2784 (.Y(n1955), 
	.A(\addr_calc/fft_read_calc/count[19] ));
   INVX2TS U2785 (.Y(n1958), 
	.A(n1957));
   INVX2TS U2787 (.Y(n1961), 
	.A(\addr_calc/iir_write_calc/count[21] ));
   INVX2TS U2788 (.Y(n1962), 
	.A(n1961));
   INVX2TS U2789 (.Y(n1963), 
	.A(\addr_calc/fft_read_calc/count[15] ));
   INVX2TS U2790 (.Y(n1965), 
	.A(n1964));
   INVX2TS U2791 (.Y(n1966), 
	.A(\addr_calc/fft_read_calc/count[13] ));
   CLKINVX3TS U2792 (.Y(n1967), 
	.A(n1966));
   INVX2TS U2793 (.Y(n1968), 
	.A(\addr_calc/iir_write_calc/count[25] ));
   INVX2TS U2794 (.Y(n1975), 
	.A(\addr_calc/fft_read_calc/count[7] ));
   INVX2TS U2796 (.Y(n1978), 
	.A(\add_x_22_0/n114 ));
   INVX2TS U2797 (.Y(n1979), 
	.A(\add_x_22_0/n121 ));
   INVX2TS U2798 (.Y(\add_x_22_0/n121 ), 
	.A(\addr_calc/fft_read_calc/count[1] ));
   NOR2X2TS U2800 (.Y(\add_x_19_1/n151 ), 
	.B(\addr_calc/fft_write_calc/count[9] ), 
	.A(FE_OFN422_offset_9_));
   INVX2TS U2803 (.Y(n1987), 
	.A(\addr_calc/fir_read_calc/count[18] ));
   INVX2TS U2804 (.Y(n1988), 
	.A(n1987));
   INVX2TS U2805 (.Y(n1991), 
	.A(\addr_calc/fir_read_calc/count[14] ));
   INVX2TS U2809 (.Y(\add_x_22_2/n101 ), 
	.A(\addr_calc/fir_read_calc/count[6] ));
   INVX2TS U2810 (.Y(n2003), 
	.A(n2002));
   INVX2TS U2811 (.Y(n2004), 
	.A(\add_x_22_2/n117 ));
   INVX2TS U2812 (.Y(\add_x_22_2/n117 ), 
	.A(\addr_calc/fir_read_calc/count[2] ));
   INVX2TS U2813 (.Y(n2810), 
	.A(\addr_calc/fir_read_calc/count[0] ));
   INVX2TS U2817 (.Y(n2012), 
	.A(\addr_calc/fir_write_calc/count[22] ));
   INVX2TS U2819 (.Y(n2015), 
	.A(\add_x_22_4/n117 ));
   INVX2TS U2820 (.Y(\add_x_22_4/n117 ), 
	.A(\addr_calc/iir_read_calc/count[2] ));
   INVX2TS U2822 (.Y(\add_x_22_4/n101 ), 
	.A(\addr_calc/iir_read_calc/count[6] ));
   INVX2TS U2823 (.Y(n2019), 
	.A(\addr_calc/fft_write_calc/count[18] ));
   AO22X1TS U2825 (.Y(n1052), 
	.B1(FE_OFN258_addr_calc_fft_write_calc_count_14_), 
	.B0(FE_OFN18_n2797), 
	.A1(\addr_calc/fft_write_calc/counter/N57 ), 
	.A0(FE_OFN27_n2795));
   NAND2X1TS U2826 (.Y(\add_x_19_1/n155 ), 
	.B(FE_OFN427_offset_8_), 
	.A(\addr_calc/fft_write_calc/count[8] ));
   INVX2TS U2827 (.Y(n2027), 
	.A(\addr_calc/iir_read_calc/count[20] ));
   NOR2X6TS U2829 (.Y(\add_x_19_4/n81 ), 
	.B(\addr_calc/iir_read_calc/count[22] ), 
	.A(FE_OCPUNCON1877_FE_OFN374_offset_22_));
   INVX2TS U2830 (.Y(n2032), 
	.A(\add_x_22_1/n117 ));
   INVX2TS U2831 (.Y(\add_x_22_1/n117 ), 
	.A(\addr_calc/fft_write_calc/count[2] ));
   INVX2TS U2832 (.Y(n2033), 
	.A(\addr_calc/iir_read_calc/count[24] ));
   INVX2TS U2833 (.Y(n2034), 
	.A(n2033));
   INVX2TS U2834 (.Y(n2036), 
	.A(\add_x_22_5/n117 ));
   INVX2TS U2835 (.Y(\add_x_22_5/n117 ), 
	.A(\addr_calc/iir_write_calc/count[2] ));
   INVX2TS U2836 (.Y(n2037), 
	.A(\addr_calc/fft_read_calc/count[24] ));
   CLKINVX3TS U2837 (.Y(n2038), 
	.A(n2037));
   INVX2TS U2838 (.Y(\add_x_22_5/n101 ), 
	.A(\addr_calc/iir_write_calc/count[6] ));
   INVX2TS U2839 (.Y(n2042), 
	.A(\addr_calc/fft_read_calc/count[14] ));
   INVX2TS U2840 (.Y(\add_x_22_5/n74 ), 
	.A(\addr_calc/iir_write_calc/count[12] ));
   INVX2TS U2841 (.Y(n2045), 
	.A(\addr_calc/fft_read_calc/count[12] ));
   INVX2TS U2842 (.Y(n2051), 
	.A(n2050));
   INVX2TS U2844 (.Y(n2056), 
	.A(\add_x_22_0/n117 ));
   INVX2TS U2845 (.Y(\add_x_22_0/n117 ), 
	.A(\addr_calc/fft_read_calc/count[2] ));
   INVX2TS U2846 (.Y(\DP_OP_158_296_6262/n1875 ), 
	.A(FE_OFN112_DP_OP_158_296_6262_n1791));
   INVX6TS U2848 (.Y(iir_enable), 
	.A(n2062));
   INVX2TS U2850 (.Y(n2071), 
	.A(FE_OFN567_n2070));
   INVX2TS U2851 (.Y(n2073), 
	.A(FE_OFN567_n2070));
   INVXLTS U2861 (.Y(n2093), 
	.A(instruction[18]));
   INVXLTS U2869 (.Y(n2108), 
	.A(instruction[19]));
   INVX2TS U2970 (.Y(n2341), 
	.A(\DP_OP_158_296_6262/n1830 ));
   INVXLTS U2972 (.Y(n2311), 
	.A(instruction[1]));
   CLKINVX2TS U2979 (.Y(n2324), 
	.A(FE_OFN462_filesize_31_));
   CLKINVX2TS U2987 (.Y(\DP_OP_158_296_6262/n1830 ), 
	.A(FE_OFN463_filesize_30_));
   INVXLTS U2989 (.Y(n2345), 
	.A(data_bus[15]));
   INVX2TS U2990 (.Y(n2347), 
	.A(data_bus[19]));
   INVXLTS U2991 (.Y(n2349), 
	.A(data_bus[11]));
   INVXLTS U2992 (.Y(n2351), 
	.A(data_bus[23]));
   INVXLTS U2993 (.Y(n2353), 
	.A(data_bus[7]));
   INVXLTS U2994 (.Y(n2355), 
	.A(data_bus[27]));
   INVXLTS U2995 (.Y(n2357), 
	.A(data_bus[3]));
   INVXLTS U2996 (.Y(n2359), 
	.A(data_bus[31]));
   INVXLTS U2997 (.Y(\DP_OP_159_297_3515/n873 ), 
	.A(FE_OFN489_filesize_11_));
   INVXLTS U2998 (.Y(\DP_OP_159_297_3515/n879 ), 
	.A(FE_OFN495_filesize_5_));
   INVXLTS U3000 (.Y(\DP_OP_159_297_3515/n877 ), 
	.A(FE_OFN493_filesize_7_));
   NOR2XLTS U3001 (.Y(\DP_OP_159_297_3515/n1069 ), 
	.B(FE_OCPUNCON1058_filesize_3_), 
	.A(\DP_OP_159_297_3515/n1074 ));
   INVXLTS U3002 (.Y(\DP_OP_159_297_3515/n867 ), 
	.A(FE_OFN480_filesize_17_));
   INVXLTS U3003 (.Y(\DP_OP_159_297_3515/n815 ), 
	.A(FE_OFN502_filesize_0_));
   INVXLTS U3039 (.Y(n2501), 
	.A(data_bus[30]));
   INVXLTS U3040 (.Y(n2503), 
	.A(data_bus[26]));
   INVXLTS U3041 (.Y(n2505), 
	.A(data_bus[22]));
   INVXLTS U3042 (.Y(n2507), 
	.A(data_bus[18]));
   INVXLTS U3043 (.Y(n2509), 
	.A(data_bus[14]));
   INVXLTS U3044 (.Y(n2511), 
	.A(data_bus[10]));
   INVXLTS U3045 (.Y(n2513), 
	.A(data_bus[6]));
   INVXLTS U3046 (.Y(n2515), 
	.A(data_bus[2]));
   INVXLTS U3047 (.Y(n2517), 
	.A(data_bus[29]));
   INVXLTS U3048 (.Y(n2519), 
	.A(data_bus[25]));
   INVXLTS U3049 (.Y(n2521), 
	.A(data_bus[21]));
   INVXLTS U3050 (.Y(n2523), 
	.A(data_bus[17]));
   INVX2TS U3051 (.Y(n2525), 
	.A(data_bus[13]));
   INVXLTS U3052 (.Y(n2527), 
	.A(data_bus[9]));
   INVXLTS U3053 (.Y(n2529), 
	.A(data_bus[5]));
   INVXLTS U3054 (.Y(n2531), 
	.A(data_bus[1]));
   INVXLTS U3055 (.Y(n2533), 
	.A(data_bus[28]));
   INVXLTS U3056 (.Y(n2535), 
	.A(data_bus[24]));
   INVXLTS U3057 (.Y(n2537), 
	.A(data_bus[20]));
   INVXLTS U3058 (.Y(n2539), 
	.A(data_bus[16]));
   INVXLTS U3059 (.Y(n2541), 
	.A(data_bus[12]));
   INVXLTS U3060 (.Y(n2543), 
	.A(data_bus[8]));
   INVXLTS U3061 (.Y(n2545), 
	.A(data_bus[4]));
   INVXLTS U3062 (.Y(n2547), 
	.A(data_bus[0]));
   NOR2X2TS U3065 (.Y(\add_x_19_0/n175 ), 
	.B(FE_OFN264_addr_calc_fft_read_calc_count_4_), 
	.A(FE_OCPUNCON1425_FE_OFN443_offset_4_));
   INVX2TS U3066 (.Y(n2554), 
	.A(\add_x_22_0/n57 ));
   NOR2X1TS U3067 (.Y(\add_x_19_0/n110 ), 
	.B(FE_OFN396_offset_16_), 
	.A(\addr_calc/fft_read_calc/count[16] ));
   INVX2TS U3068 (.Y(n2555), 
	.A(\add_x_22_1/n30 ));
   INVX2TS U3069 (.Y(n2556), 
	.A(\add_x_22_4/n46 ));
   INVX2TS U3070 (.Y(n2557), 
	.A(\add_x_22_1/n7 ));
   INVX2TS U3071 (.Y(n2558), 
	.A(\add_x_22_2/n30 ));
   NOR2X1TS U3072 (.Y(\add_x_19_2/n78 ), 
	.B(FE_OFN369_offset_23_), 
	.A(\addr_calc/fir_read_calc/count[23] ));
   INVX2TS U3073 (.Y(n2559), 
	.A(\add_x_22_0/n7 ));
   INVX2TS U3074 (.Y(n2560), 
	.A(\add_x_22_0/n89 ));
   INVX2TS U3075 (.Y(n2561), 
	.A(\add_x_22_4/n7 ));
   INVX2TS U3076 (.Y(n2562), 
	.A(\add_x_22_5/n89 ));
   INVX2TS U3077 (.Y(n2563), 
	.A(\add_x_22_3/n30 ));
   INVX2TS U3078 (.Y(n2564), 
	.A(\add_x_22_3/n57 ));
   NAND2X1TS U3079 (.Y(\add_x_19_3/n111 ), 
	.B(FE_OFN396_offset_16_), 
	.A(\addr_calc/fir_write_calc/count[16] ));
   INVX2TS U3080 (.Y(n2565), 
	.A(\add_x_22_4/n30 ));
   INVX2TS U3081 (.Y(n2567), 
	.A(\add_x_22_1/n57 ));
   NAND2X1TS U3082 (.Y(\add_x_19_1/n111 ), 
	.B(\addr_calc/fft_write_calc/count[16] ), 
	.A(FE_OFN395_offset_16_));
   INVX2TS U3083 (.Y(n2568), 
	.A(\add_x_22_1/n114 ));
   INVX2TS U3084 (.Y(n2570), 
	.A(\add_x_22_5/n67 ));
   INVX2TS U3086 (.Y(n2572), 
	.A(\add_x_22_0/n40 ));
   INVX2TS U3087 (.Y(n2573), 
	.A(\add_x_22_5/n15 ));
   INVX2TS U3088 (.Y(n2574), 
	.A(\add_x_22_1/n15 ));
   INVX2TS U3089 (.Y(n2575), 
	.A(\add_x_22_0/n15 ));
   INVX2TS U3091 (.Y(n2577), 
	.A(\add_x_22_3/n22 ));
   INVX2TS U3092 (.Y(n2578), 
	.A(n2791));
   XNOR2X1TS U3093 (.Y(\DP_OP_159_297_3515/n778 ), 
	.B(\DP_OP_159_297_3515/n815 ), 
	.A(\addr_calc/iir_write_calc/count[0] ));
   INVX2TS U3094 (.Y(n2579), 
	.A(\add_x_22_5/n33 ));
   INVX2TS U3095 (.Y(n2580), 
	.A(n2786));
   NOR4X1TS U3097 (.Y(n863), 
	.D(\addr_calc/fir_write_calc/count[24] ), 
	.C(n1835), 
	.B(FE_OFN267_addr_calc_fir_write_calc_count_26_), 
	.A(FE_OFN231_addr_calc_fir_write_calc_count_25_));
   NOR2X1TS U3099 (.Y(\add_x_19_2/n58 ), 
	.B(FE_OFN357_offset_26_), 
	.A(FE_OFN269_addr_calc_fir_read_calc_count_26_));
   INVX2TS U3100 (.Y(n2583), 
	.A(\add_x_22_4/n92 ));
   INVX2TS U3101 (.Y(n2587), 
	.A(FE_OFN151_n2074));
   AOI211XLTS U3103 (.Y(\data_cntl/N252 ), 
	.C0(n2587), 
	.B0(FE_OFN507_from_fft_empty), 
	.A1(n938), 
	.A0(FE_OFN505_to_fft_empty));
   INVX2TS U3104 (.Y(\add_x_22_0/n57 ), 
	.A(\addr_calc/fft_read_calc/count[16] ));
   INVX2TS U3105 (.Y(\add_x_22_0/n23 ), 
	.A(\add_x_22_0/n24 ));
   XNOR2X1TS U3106 (.Y(\addr_calc/fir_read_calc/counter/N44 ), 
	.B(n2007), 
	.A(\add_x_22_2/n121 ));
   INVX2TS U3108 (.Y(\add_x_22_2/n30 ), 
	.A(\addr_calc/fir_read_calc/count[23] ));
   INVX2TS U3110 (.Y(\add_x_22_3/n57 ), 
	.A(\addr_calc/fir_write_calc/count[16] ));
   INVX2TS U3111 (.Y(\add_x_22_3/n22 ), 
	.A(\addr_calc/fir_write_calc/count[24] ));
   INVX2TS U3112 (.Y(\add_x_22_5/n53 ), 
	.A(\addr_calc/iir_write_calc/count[17] ));
   INVX2TS U3113 (.Y(\add_x_22_5/n33 ), 
	.A(\addr_calc/iir_write_calc/count[22] ));
   INVX2TS U3114 (.Y(\add_x_22_1/n57 ), 
	.A(\addr_calc/fft_write_calc/count[16] ));
   INVX2TS U3115 (.Y(\add_x_22_4/n33 ), 
	.A(\addr_calc/iir_read_calc/count[22] ));
   INVX2TS U3116 (.Y(\add_x_22_4/n57 ), 
	.A(\addr_calc/iir_read_calc/count[16] ));
   INVXLTS U3117 (.Y(\add_x_22_4/n105 ), 
	.A(\addr_calc/iir_read_calc/count[5] ));
   XNOR2X1TS U3118 (.Y(\DP_OP_158_296_6262/n375 ), 
	.B(\addr_calc/fir_read_calc/count[0] ), 
	.A(FE_OFN518_n2372));
   XOR2X1TS U3119 (.Y(n2590), 
	.B(n2004), 
	.A(n2596));
   XOR2X1TS U3120 (.Y(n2591), 
	.B(\addr_calc/fir_read_calc/count[6] ), 
	.A(n2593));
   XOR2X1TS U3121 (.Y(n2592), 
	.B(n1908), 
	.A(FE_OFN75_n2599));
   XOR2X1TS U3122 (.Y(n2600), 
	.B(\addr_calc/fir_read_calc/count[4] ), 
	.A(\DP_OP_158_296_6262/n855 ));
   XOR2X1TS U3123 (.Y(n2601), 
	.B(FE_OFN245_addr_calc_fir_read_calc_count_5_), 
	.A(n2595));
   INVXLTS U3124 (.Y(\DP_OP_158_296_6262/n1972 ), 
	.A(n1138));
   CLKXOR2X2TS U3125 (.Y(n2597), 
	.B(FE_OFN502_filesize_0_), 
	.A(FE_OFN501_filesize_1_));
   INVX2TS U3126 (.Y(\DP_OP_158_296_6262/n2010 ), 
	.A(\DP_OP_158_296_6262/n2011 ));
   CLKINVX4TS U3127 (.Y(\DP_OP_158_296_6262/n855 ), 
	.A(\DP_OP_158_296_6262/n2034 ));
   INVXLTS U3128 (.Y(\DP_OP_158_296_6262/n1863 ), 
	.A(\DP_OP_158_296_6262/n1862 ));
   INVXLTS U3129 (.Y(\DP_OP_158_296_6262/n1917 ), 
	.A(\DP_OP_158_296_6262/n1918 ));
   INVX2TS U3130 (.Y(\DP_OP_158_296_6262/n2020 ), 
	.A(n1797));
   CLKINVX2TS U3131 (.Y(\DP_OP_158_296_6262/n1904 ), 
	.A(\DP_OP_158_296_6262/n1903 ));
   CLKINVX2TS U3132 (.Y(\DP_OP_158_296_6262/n1849 ), 
	.A(\DP_OP_158_296_6262/n1792 ));
   XOR2X4TS U3133 (.Y(\DP_OP_158_296_6262/n2054 ), 
	.B(FE_OFN471_filesize_24_), 
	.A(\DP_OP_158_296_6262/n1874 ));
   NOR2X2TS U3134 (.Y(\DP_OP_158_296_6262/n66 ), 
	.B(\DP_OP_158_296_6262/n87 ), 
	.A(\DP_OP_158_296_6262/n68 ));
   NOR2X4TS U3135 (.Y(\DP_OP_158_296_6262/n3 ), 
	.B(\DP_OP_158_296_6262/n5 ), 
	.A(\DP_OP_158_296_6262/n18 ));
   NOR2X2TS U3136 (.Y(\DP_OP_158_296_6262/n37 ), 
	.B(\DP_OP_158_296_6262/n39 ), 
	.A(\DP_OP_158_296_6262/n54 ));
   NOR2X1TS U3137 (.Y(\DP_OP_158_296_6262/n159 ), 
	.B(\DP_OP_158_296_6262/n161 ), 
	.A(\DP_OP_158_296_6262/n174 ));
   NAND2X1TS U3138 (.Y(\DP_OP_159_297_3515/n892 ), 
	.B(\DP_OP_159_297_3515/n893 ), 
	.A(FE_OCPUNCON1566_n1789));
   XOR2X1TS U3139 (.Y(n2604), 
	.B(\addr_calc/iir_write_calc/count[2] ), 
	.A(n2612));
   XOR2X1TS U3140 (.Y(n2605), 
	.B(n2039), 
	.A(n2610));
   XOR2X1TS U3141 (.Y(n2606), 
	.B(n1935), 
	.A(n2624));
   XOR2X1TS U3142 (.Y(n2609), 
	.B(\DP_OP_159_297_3515/n877 ), 
	.A(\DP_OP_159_297_3515/n1051 ));
   XOR2X1TS U3143 (.Y(n2611), 
	.B(FE_OCPUNCON1058_filesize_3_), 
	.A(\DP_OP_159_297_3515/n1074 ));
   XOR2X1TS U3144 (.Y(n2612), 
	.B(FE_OFN500_filesize_1_), 
	.A(n1680));
   XNOR2X1TS U3145 (.Y(n2623), 
	.B(\DP_OP_159_297_3515/n879 ), 
	.A(\DP_OP_159_297_3515/n1063 ));
   XNOR2X1TS U3146 (.Y(n2624), 
	.B(\DP_OP_159_297_3515/n880 ), 
	.A(\DP_OP_159_297_3515/n1069 ));
   XOR2X1TS U3147 (.Y(n2626), 
	.B(n1686), 
	.A(n2623));
   INVX2TS U3148 (.Y(\DP_OP_159_297_3515/n1012 ), 
	.A(\DP_OP_159_297_3515/n1011 ));
   INVX2TS U3149 (.Y(\DP_OP_159_297_3515/n1063 ), 
	.A(\DP_OP_159_297_3515/n1064 ));
   INVXLTS U3150 (.Y(\DP_OP_159_297_3515/n1074 ), 
	.A(\DP_OP_159_297_3515/n1075 ));
   INVXLTS U3151 (.Y(\DP_OP_159_297_3515/n916 ), 
	.A(\DP_OP_159_297_3515/n915 ));
   INVXLTS U3152 (.Y(\DP_OP_159_297_3515/n999 ), 
	.A(\DP_OP_159_297_3515/n998 ));
   XOR2X4TS U3153 (.Y(\DP_OP_159_297_3515/n1138 ), 
	.B(n2330), 
	.A(\DP_OP_159_297_3515/n906 ));
   NOR2X1TS U3154 (.Y(\DP_OP_159_297_3515/n740 ), 
	.B(\DP_OP_159_297_3515/n758 ), 
	.A(\DP_OP_159_297_3515/n742 ));
   NAND2X1TS U3155 (.Y(\DP_OP_159_297_3515/n726 ), 
	.B(\DP_OP_159_297_3515/n740 ), 
	.A(\DP_OP_159_297_3515/n728 ));
   XNOR2X1TS U3156 (.Y(\DP_OP_159_297_3515/n610 ), 
	.B(\addr_calc/iir_write_calc/count[19] ), 
	.A(n1662));
   OR2X2TS U3157 (.Y(n2628), 
	.B(FE_OFN348_offset_29_), 
	.A(FE_OFN275_addr_calc_fft_read_calc_count_29_));
   OR2X2TS U3158 (.Y(n2627), 
	.B(FE_OFN339_offset_31_), 
	.A(FE_OFN226_addr_calc_fft_read_calc_count_31_));
   CLKINVX8TS U3159 (.Y(\add_x_19_0/n68 ), 
	.A(\add_x_19_0/n69 ));
   CLKINVX20TS U3163 (.Y(\add_x_19_5/n156 ), 
	.A(FE_OFN129_add_x_19_5_n157));
   OR2X2TS U3164 (.Y(n2629), 
	.B(FE_OFN347_offset_29_), 
	.A(n1851));
   INVX6TS U3165 (.Y(\add_x_19_5/n112 ), 
	.A(\add_x_19_5/n113 ));
   CLKINVX3TS U3166 (.Y(\add_x_19_5/n91 ), 
	.A(\add_x_19_5/n92 ));
   INVX6TS U3167 (.Y(\add_x_19_5/n68 ), 
	.A(\add_x_19_5/n69 ));
   INVX12TS U3170 (.Y(\add_x_19_3/n156 ), 
	.A(FE_OFN525_add_x_19_3_n157));
   OR2X2TS U3171 (.Y(n2631), 
	.B(FE_OFN348_offset_29_), 
	.A(FE_OFN273_addr_calc_fir_write_calc_count_29_));
   AOI21X4TS U3173 (.Y(\add_x_19_3/n60 ), 
	.B0(\add_x_19_3/n62 ), 
	.A1(\add_x_19_3/n61 ), 
	.A0(\add_x_19_3/n69 ));
   INVXLTS U3174 (.Y(\add_x_19_1/n212 ), 
	.A(\add_x_19_1/n139 ));
   OR2X2TS U3175 (.Y(n2632), 
	.B(FE_OFN345_offset_29_), 
	.A(\addr_calc/fft_write_calc/count[29] ));
   OR2XLTS U3176 (.Y(n2633), 
	.B(FE_OFN346_offset_29_), 
	.A(n1842));
   INVX4TS U3177 (.Y(\add_x_19_2/n68 ), 
	.A(\add_x_19_2/n69 ));
   OR2X2TS U3179 (.Y(n2634), 
	.B(FE_OFN347_offset_29_), 
	.A(\addr_calc/iir_read_calc/count[29] ));
   INVX4TS U3180 (.Y(\add_x_19_4/n133 ), 
	.A(\add_x_19_4/n134 ));
   AO22X1TS U3182 (.Y(n972), 
	.B1(\addr_calc/iir_read_calc/count[31] ), 
	.B0(FE_OFN89_n2654), 
	.A1(\addr_calc/iir_read_calc/counter/N74 ), 
	.A0(FE_OFN82_n2787));
   AO22X1TS U3183 (.Y(n988), 
	.B1(n2570), 
	.B0(FE_OCPUNCON1569_n2812), 
	.A1(\addr_calc/iir_write_calc/counter/N57 ), 
	.A0(FE_OCPUNCON1881_n2813));
   AO22X1TS U3184 (.Y(n941), 
	.B1(\addr_calc/iir_read_calc/count[30] ), 
	.B0(FE_OFN92_n1192), 
	.A1(\addr_calc/iir_read_calc/counter/N73 ), 
	.A0(FE_OFN82_n2787));
   AO22X4TS U3185 (.Y(n995), 
	.B1(n1683), 
	.B0(FE_OCPUNCON1576_n2812), 
	.A1(\addr_calc/iir_write_calc/counter/N50 ), 
	.A0(FE_OCPUNCON1888_n2813));
   AO22X1TS U3186 (.Y(n990), 
	.B1(n2044), 
	.B0(FE_OCPUNCON1569_n2812), 
	.A1(\addr_calc/iir_write_calc/counter/N55 ), 
	.A0(FE_OCPUNCON1879_n2813));
   AO22X1TS U3187 (.Y(n992), 
	.B1(n1940), 
	.B0(n2812), 
	.A1(\addr_calc/iir_write_calc/counter/N53 ), 
	.A0(n2813));
   AO22X1TS U3188 (.Y(n973), 
	.B1(n1851), 
	.B0(FE_OCPUNCON1574_n2812), 
	.A1(\addr_calc/iir_write_calc/counter/N72 ), 
	.A0(FE_OCPUNCON1885_n2813));
   AO22X1TS U3189 (.Y(n961), 
	.B1(\addr_calc/iir_read_calc/count[10] ), 
	.B0(n1192), 
	.A1(\addr_calc/iir_read_calc/counter/N53 ), 
	.A0(n2787));
   AO22X1TS U3190 (.Y(n963), 
	.B1(n2583), 
	.B0(FE_OFN85_n2654), 
	.A1(\addr_calc/iir_read_calc/counter/N51 ), 
	.A0(n2787));
   AO22X1TS U3191 (.Y(n962), 
	.B1(n1685), 
	.B0(n2654), 
	.A1(\addr_calc/iir_read_calc/counter/N52 ), 
	.A0(FE_OCPUNCON1878_n2787));
   CLKINVX2TS U3193 (.Y(n785), 
	.A(\addr_calc/fir_write_calc/counter/N38 ));
   AO22X1TS U3194 (.Y(n956), 
	.B1(n2566), 
	.B0(FE_OFN90_n1192), 
	.A1(\addr_calc/iir_read_calc/counter/N58 ), 
	.A0(FE_OCPUNCON1880_n2787));
   NOR4X1TS U3195 (.Y(n878), 
	.D(n1983), 
	.C(n1876), 
	.B(FE_OFN270_addr_calc_fir_read_calc_count_26_), 
	.A(FE_OFN243_addr_calc_fir_read_calc_count_27_));
   NOR4X1TS U3196 (.Y(n876), 
	.D(FE_OFN261_addr_calc_fir_read_calc_count_31_), 
	.C(n1908), 
	.B(n1906), 
	.A(FE_OFN245_addr_calc_fir_read_calc_count_5_));
   NOR4X1TS U3197 (.Y(n861), 
	.D(FE_OFN262_addr_calc_fir_write_calc_count_31_), 
	.C(n1866), 
	.B(FE_OFN241_addr_calc_fir_write_calc_count_4_), 
	.A(n1867));
   NOR4XLTS U3198 (.Y(n831), 
	.D(\addr_calc/fft_read_calc/count[28] ), 
	.C(FE_OFN275_addr_calc_fft_read_calc_count_29_), 
	.B(n2056), 
	.A(FE_OFN278_addr_calc_fft_read_calc_count_30_));
   NOR4X1TS U3199 (.Y(n830), 
	.D(n2038), 
	.C(\addr_calc/fft_read_calc/count[25] ), 
	.B(\addr_calc/fft_read_calc/count[26] ), 
	.A(\addr_calc/fft_read_calc/count[27] ));
   NOR4X1TS U3200 (.Y(n828), 
	.D(FE_OFN226_addr_calc_fft_read_calc_count_31_), 
	.C(n1978), 
	.B(FE_OFN263_addr_calc_fft_read_calc_count_4_), 
	.A(FE_OFN251_addr_calc_fft_read_calc_count_5_));
   NOR4X1TS U3201 (.Y(n845), 
	.D(\addr_calc/fft_write_calc/count[28] ), 
	.C(n1853), 
	.B(n2032), 
	.A(FE_OFN279_addr_calc_fft_write_calc_count_30_));
   NOR4X1TS U3202 (.Y(n844), 
	.D(FE_OFN277_addr_calc_fft_write_calc_count_24_), 
	.C(\addr_calc/fft_write_calc/count[25] ), 
	.B(\addr_calc/fft_write_calc/count[26] ), 
	.A(\addr_calc/fft_write_calc/count[27] ));
   NOR4X2TS U3203 (.Y(n842), 
	.D(FE_OFN274_addr_calc_fft_write_calc_count_31_), 
	.C(n2568), 
	.B(n1939), 
	.A(n1479));
   NOR4X1TS U3204 (.Y(n917), 
	.D(\addr_calc/iir_write_calc/count[24] ), 
	.C(\addr_calc/iir_write_calc/count[25] ), 
	.B(\addr_calc/iir_write_calc/count[26] ), 
	.A(\addr_calc/iir_write_calc/count[27] ));
   NOR4X1TS U3206 (.Y(n813), 
	.D(\addr_calc/iir_read_calc/count[28] ), 
	.C(n1840), 
	.B(n2015), 
	.A(FE_OFN286_addr_calc_iir_read_calc_count_30_));
   NOR4X1TS U3207 (.Y(n812), 
	.D(n2034), 
	.C(\addr_calc/iir_read_calc/count[25] ), 
	.B(\addr_calc/iir_read_calc/count[26] ), 
	.A(FE_OFN235_addr_calc_iir_read_calc_count_27_));
   NOR4X1TS U3209 (.Y(n810), 
	.D(FE_OFN234_addr_calc_iir_read_calc_count_31_), 
	.C(\addr_calc/iir_read_calc/count[3] ), 
	.B(\addr_calc/iir_read_calc/count[4] ), 
	.A(n2553));
   NOR4X2TS U3210 (.Y(n915), 
	.D(FE_OFN240_addr_calc_iir_write_calc_count_31_), 
	.C(FE_OFN250_addr_calc_iir_write_calc_count_3_), 
	.B(n1935), 
	.A(\addr_calc/iir_write_calc/count[5] ));
   NOR2X1TS U3211 (.Y(n2808), 
	.B(n2799), 
	.A(n2800));
   NOR2X2TS U3212 (.Y(n2804), 
	.B(n2801), 
	.A(n2802));
   NOR2X1TS U3213 (.Y(n2785), 
	.B(n2783), 
	.A(n2784));
   AO22X1TS U3217 (.Y(n1079), 
	.B1(n1881), 
	.B0(FE_OFN65_n2809), 
	.A1(\addr_calc/fir_read_calc/counter/N62 ), 
	.A0(FE_OFN55_n2807));
   AO22X2TS U3218 (.Y(n1101), 
	.B1(\addr_calc/fir_write_calc/count[29] ), 
	.B0(FE_OCPUNCON1090_n2805), 
	.A1(\addr_calc/fir_write_calc/counter/N72 ), 
	.A0(n1762));
   AO22X1TS U3219 (.Y(n1019), 
	.B1(n1689), 
	.B0(FE_OFN7_n2794), 
	.A1(\addr_calc/fft_read_calc/counter/N58 ), 
	.A0(n1755));
   AO22X2TS U3220 (.Y(n1005), 
	.B1(\addr_calc/fft_read_calc/count[29] ), 
	.B0(FE_OFN14_n2794), 
	.A1(\addr_calc/fft_read_calc/counter/N72 ), 
	.A0(FE_OFN4_n1755));
   AO22X2TS U3221 (.Y(n1037), 
	.B1(n1853), 
	.B0(FE_OFN24_n2797), 
	.A1(\addr_calc/fft_write_calc/counter/N72 ), 
	.A0(FE_OFN33_n2795));
   INVX2TS U3226 (.Y(n451), 
	.A(FE_OFN314_data_cntl_N159));
   INVX2TS U3240 (.Y(n643), 
	.A(FE_OFN332_data_cntl_N63));
   INVX2TS U3246 (.Y(n515), 
	.A(FE_OFN329_data_cntl_N99));
   INVX2TS U3252 (.Y(n387), 
	.A(FE_OFN326_data_cntl_N191));
   INVX2TS U3257 (.Y(n707), 
	.A(FE_OFN322_data_cntl_N9));
   INVX2TS U3262 (.Y(n579), 
	.A(FE_OFN318_data_cntl_N95));
   INVX2TS U3266 (.Y(n131), 
	.A(\addr_calc/N99 ));
   INVX2TS U3272 (.Y(n195), 
	.A(\addr_calc/N95 ));
   INVX2TS U3275 (.Y(n259), 
	.A(\addr_calc/N63 ));
   INVX2TS U3279 (.Y(n323), 
	.A(\addr_calc/N9 ));
   INVX2TS U3281 (.Y(n67), 
	.A(\addr_calc/N159 ));
   INVX2TS U3284 (.Y(n3), 
	.A(\addr_calc/N191 ));
   AO22X1TS U3285 (.Y(n1096), 
	.B1(n2004), 
	.B0(FE_OFN70_n2809), 
	.A1(\addr_calc/fir_read_calc/counter/N45 ), 
	.A0(FE_OFN60_n2807));
   AO22X1TS U3286 (.Y(n1086), 
	.B1(n1994), 
	.B0(FE_OFN62_n2809), 
	.A1(\addr_calc/fir_read_calc/counter/N55 ), 
	.A0(FE_OFN52_n2807));
   AO22X2TS U3287 (.Y(n1092), 
	.B1(n2001), 
	.B0(FE_OFN71_n2809), 
	.A1(\addr_calc/fir_read_calc/counter/N49 ), 
	.A0(FE_OFN61_n2807));
   AO22X1TS U3288 (.Y(n1081), 
	.B1(n1884), 
	.B0(FE_OFN65_n2809), 
	.A1(\addr_calc/fir_read_calc/counter/N60 ), 
	.A0(FE_OFN55_n2807));
   AO22X1TS U3289 (.Y(n1085), 
	.B1(n1893), 
	.B0(n2809), 
	.A1(\addr_calc/fir_read_calc/counter/N56 ), 
	.A0(FE_OFN52_n2807));
   AO22X1TS U3290 (.Y(n1087), 
	.B1(n1895), 
	.B0(FE_OFN62_n2809), 
	.A1(\addr_calc/fir_read_calc/counter/N54 ), 
	.A0(n2807));
   AO22X1TS U3291 (.Y(n1090), 
	.B1(n1997), 
	.B0(FE_OFN63_n2809), 
	.A1(\addr_calc/fir_read_calc/counter/N51 ), 
	.A0(FE_OFN54_n2807));
   AO22X1TS U3292 (.Y(n1074), 
	.B1(\addr_calc/fir_read_calc/count[24] ), 
	.B0(FE_OFN68_n2809), 
	.A1(\addr_calc/fir_read_calc/counter/N67 ), 
	.A0(FE_OFN58_n2807));
   AO22X2TS U3293 (.Y(n1127), 
	.B1(n1866), 
	.B0(FE_OCPUNCON1091_n2805), 
	.A1(\addr_calc/fir_write_calc/counter/N46 ), 
	.A0(FE_OFN549_n1763));
   AO22X1TS U3294 (.Y(n1122), 
	.B1(FE_OFN256_addr_calc_fir_write_calc_count_8_), 
	.B0(n2805), 
	.A1(\addr_calc/fir_write_calc/counter/N51 ), 
	.A0(FE_OFN547_n2803));
   AO22X1TS U3295 (.Y(n1119), 
	.B1(n1877), 
	.B0(FE_OCPUNCON1083_n2805), 
	.A1(\addr_calc/fir_write_calc/counter/N54 ), 
	.A0(FE_OFN547_n2803));
   AO22X2TS U3297 (.Y(n1124), 
	.B1(FE_OFN253_addr_calc_fir_write_calc_count_6_), 
	.B0(FE_OCPUNCON1092_n2805), 
	.A1(\addr_calc/fir_write_calc/counter/N49 ), 
	.A0(FE_OFN51_n2803));
   AO22X1TS U3298 (.Y(n1117), 
	.B1(n1880), 
	.B0(FE_OCPUNCON1083_n2805), 
	.A1(\addr_calc/fir_write_calc/counter/N56 ), 
	.A0(FE_OFN548_n1763));
   AO22X1TS U3299 (.Y(n1103), 
	.B1(\addr_calc/fir_write_calc/count[27] ), 
	.B0(FE_OCPUNCON1089_n2805), 
	.A1(\addr_calc/fir_write_calc/counter/N70 ), 
	.A0(FE_OFN50_n2803));
   AO22X1TS U3300 (.Y(n1107), 
	.B1(n2563), 
	.B0(FE_OCPUNCON1086_n2805), 
	.A1(\addr_calc/fir_write_calc/counter/N66 ), 
	.A0(FE_OFN49_n2803));
   AO22X1TS U3301 (.Y(n1102), 
	.B1(n1896), 
	.B0(FE_OCPUNCON1088_n2805), 
	.A1(\addr_calc/fir_write_calc/counter/N71 ), 
	.A0(FE_OFN549_n1763));
   AO22X1TS U3302 (.Y(n1099), 
	.B1(\addr_calc/fir_write_calc/count[31] ), 
	.B0(FE_OCPUNCON1090_n2805), 
	.A1(\addr_calc/fir_write_calc/counter/N74 ), 
	.A0(FE_OFN51_n2803));
   AO22X2TS U3303 (.Y(n1033), 
	.B1(FE_OFN16_n2794), 
	.B0(n1979), 
	.A1(\addr_calc/fft_read_calc/counter/N44 ), 
	.A0(FE_OFN3_n1754));
   AO22X2TS U3304 (.Y(n1032), 
	.B1(FE_OFN16_n2794), 
	.B0(n2056), 
	.A1(\addr_calc/fft_read_calc/counter/N45 ), 
	.A0(FE_OFN3_n1754));
   AO22X1TS U3305 (.Y(n1114), 
	.B1(n2564), 
	.B0(FE_OCPUNCON1085_n2805), 
	.A1(\addr_calc/fir_write_calc/counter/N59 ), 
	.A0(FE_OFN48_n2803));
   AO22X1TS U3306 (.Y(n1106), 
	.B1(n2577), 
	.B0(FE_OCPUNCON1088_n2805), 
	.A1(\addr_calc/fir_write_calc/counter/N67 ), 
	.A0(FE_OFN50_n2803));
   AO22X1TS U3307 (.Y(n1113), 
	.B1(FE_OCPUNCON1085_n2805), 
	.B0(\addr_calc/fir_write_calc/count[17] ), 
	.A1(\addr_calc/fir_write_calc/counter/N60 ), 
	.A0(FE_OFN48_n2803));
   AO22X2TS U3308 (.Y(n1031), 
	.B1(n1978), 
	.B0(FE_OFN16_n2794), 
	.A1(\addr_calc/fft_read_calc/counter/N46 ), 
	.A0(FE_OFN550_n1750));
   AO22X1TS U3309 (.Y(n1026), 
	.B1(n2049), 
	.B0(FE_OFN9_n2794), 
	.A1(\addr_calc/fft_read_calc/counter/N51 ), 
	.A0(n1754));
   AO22X1TS U3310 (.Y(n1025), 
	.B1(n2560), 
	.B0(FE_OFN8_n2794), 
	.A1(\addr_calc/fft_read_calc/counter/N52 ), 
	.A0(FE_OFN6_n1750));
   AO22X1TS U3311 (.Y(n1024), 
	.B1(n1972), 
	.B0(FE_OFN7_n2794), 
	.A1(\addr_calc/fft_read_calc/counter/N53 ), 
	.A0(FE_OFN1_n1751));
   AO22X2TS U3312 (.Y(n1029), 
	.B1(\addr_calc/fft_read_calc/count[5] ), 
	.B0(FE_OFN15_n2794), 
	.A1(\addr_calc/fft_read_calc/counter/N48 ), 
	.A0(FE_OFN4_n1755));
   AO22X1TS U3313 (.Y(n1009), 
	.B1(FE_OFN13_n2794), 
	.B0(\addr_calc/fft_read_calc/count[25] ), 
	.A1(\addr_calc/fft_read_calc/counter/N68 ), 
	.A0(n1755));
   AO22X1TS U3314 (.Y(n1007), 
	.B1(FE_OFN13_n2794), 
	.B0(\addr_calc/fft_read_calc/count[27] ), 
	.A1(\addr_calc/fft_read_calc/counter/N70 ), 
	.A0(FE_OFN3_n1754));
   AO22X1TS U3315 (.Y(n1011), 
	.B1(\addr_calc/fft_read_calc/count[23] ), 
	.B0(FE_OFN12_n2794), 
	.A1(\addr_calc/fft_read_calc/counter/N66 ), 
	.A0(FE_OFN550_n1750));
   AO22X1TS U3316 (.Y(n1010), 
	.B1(\addr_calc/fft_read_calc/count[24] ), 
	.B0(FE_OFN12_n2794), 
	.A1(\addr_calc/fft_read_calc/counter/N67 ), 
	.A0(FE_OFN550_n1750));
   AO22X1TS U3317 (.Y(n1041), 
	.B1(\addr_calc/fft_write_calc/count[25] ), 
	.B0(FE_OFN23_n2797), 
	.A1(\addr_calc/fft_write_calc/counter/N68 ), 
	.A0(FE_OFN32_n2795));
   AO22X1TS U3318 (.Y(n1015), 
	.B1(FE_OFN10_n2794), 
	.B0(n1956), 
	.A1(\addr_calc/fft_read_calc/counter/N62 ), 
	.A0(FE_OFN552_n1751));
   AO22X2TS U3319 (.Y(n1067), 
	.B1(\addr_calc/fft_write_calc/count[31] ), 
	.B0(FE_OFN24_n2797), 
	.A1(\addr_calc/fft_write_calc/counter/N74 ), 
	.A0(FE_OFN33_n2795));
   AO22XLTS U3320 (.Y(n969), 
	.B1(FE_OFN89_n2654), 
	.B0(n2015), 
	.A1(\addr_calc/iir_read_calc/counter/N45 ), 
	.A0(FE_OFN83_n2787));
   AO22X1TS U3321 (.Y(n970), 
	.B1(FE_OFN89_n2654), 
	.B0(n1898), 
	.A1(\addr_calc/iir_read_calc/counter/N44 ), 
	.A0(FE_OFN83_n2787));
   AO22X1TS U3322 (.Y(n943), 
	.B1(n2561), 
	.B0(FE_OFN88_n2654), 
	.A1(\addr_calc/iir_read_calc/counter/N71 ), 
	.A0(FE_OFN80_n2787));
   AO22X1TS U3323 (.Y(n946), 
	.B1(\addr_calc/iir_read_calc/count[25] ), 
	.B0(FE_OFN92_n1192), 
	.A1(\addr_calc/iir_read_calc/counter/N68 ), 
	.A0(FE_OFN81_n2787));
   AO22X1TS U3324 (.Y(n947), 
	.B1(FE_OFN87_n2654), 
	.B0(\addr_calc/iir_read_calc/count[24] ), 
	.A1(\addr_calc/iir_read_calc/counter/N67 ), 
	.A0(FE_OFN80_n2787));
   AO22X1TS U3325 (.Y(n942), 
	.B1(n1840), 
	.B0(FE_OFN89_n2654), 
	.A1(\addr_calc/iir_read_calc/counter/N72 ), 
	.A0(FE_OFN82_n2787));
   AO22X1TS U3326 (.Y(n955), 
	.B1(FE_OFN86_n2654), 
	.B0(\addr_calc/iir_read_calc/count[16] ), 
	.A1(\addr_calc/iir_read_calc/counter/N59 ), 
	.A0(FE_OCPUNCON1880_n2787));
   AO22X2TS U3327 (.Y(n998), 
	.B1(n1935), 
	.B0(FE_OCPUNCON1576_n2812), 
	.A1(\addr_calc/iir_write_calc/counter/N47 ), 
	.A0(FE_OCPUNCON1888_n2813));
   AO22X1TS U3328 (.Y(n976), 
	.B1(n2573), 
	.B0(FE_OCPUNCON1573_n2812), 
	.A1(\addr_calc/iir_write_calc/counter/N69 ), 
	.A0(FE_OCPUNCON1885_n2813));
   AO22X1TS U3329 (.Y(n975), 
	.B1(n1688), 
	.B0(FE_OCPUNCON1573_n2812), 
	.A1(\addr_calc/iir_write_calc/counter/N70 ), 
	.A0(FE_OCPUNCON1884_n2813));
   AO22X1TS U3330 (.Y(n977), 
	.B1(\addr_calc/iir_write_calc/count[25] ), 
	.B0(FE_OCPUNCON1574_n2812), 
	.A1(\addr_calc/iir_write_calc/counter/N68 ), 
	.A0(FE_OCPUNCON1885_n2813));
   AO22X1TS U3331 (.Y(n1003), 
	.B1(\addr_calc/iir_write_calc/count[30] ), 
	.B0(FE_OCPUNCON1574_n2812), 
	.A1(\addr_calc/iir_write_calc/counter/N73 ), 
	.A0(FE_OCPUNCON1886_n2813));
   AO22X1TS U3332 (.Y(n983), 
	.B1(\addr_calc/iir_write_calc/count[19] ), 
	.B0(FE_OCPUNCON1571_n2812), 
	.A1(\addr_calc/iir_write_calc/counter/N62 ), 
	.A0(FE_OCPUNCON1882_n2813));
   OAI21XLTS U3384 (.Y(n2811), 
	.B0(fir_enable), 
	.A1(n2808), 
	.A0(n2810));
   OAI21XLTS U3385 (.Y(n2806), 
	.B0(FE_OFN566_n2066), 
	.A1(n2804), 
	.A0(\addr_calc/fir_write_calc/counter/N43 ));
   NAND4X1TS U3386 (.Y(n2800), 
	.D(n883), 
	.C(n882), 
	.B(n881), 
	.A(n880));
   NAND4X2TS U3387 (.Y(n2801), 
	.D(n864), 
	.C(n863), 
	.B(n862), 
	.A(n861));
   NOR4XLTS U3388 (.Y(n862), 
	.D(FE_OFN254_addr_calc_fir_write_calc_count_6_), 
	.C(\addr_calc/fir_write_calc/count[7] ), 
	.B(FE_OFN257_addr_calc_fir_write_calc_count_8_), 
	.A(n1872));
   NAND4X1TS U3389 (.Y(n2802), 
	.D(n868), 
	.C(n867), 
	.B(n866), 
	.A(n865));
   NOR4XLTS U3390 (.Y(n829), 
	.D(\addr_calc/fft_read_calc/count[6] ), 
	.C(\addr_calc/fft_read_calc/count[7] ), 
	.B(n2049), 
	.A(n2560));
   NOR4XLTS U3391 (.Y(n843), 
	.D(FE_OFN272_addr_calc_fft_write_calc_count_6_), 
	.C(n1934), 
	.B(n2026), 
	.A(n1936));
   NAND4X2TS U3392 (.Y(n2783), 
	.D(n813), 
	.C(n812), 
	.B(n811), 
	.A(n810));
   NOR4XLTS U3393 (.Y(n811), 
	.D(n2018), 
	.C(FE_OFN246_addr_calc_iir_read_calc_count_7_), 
	.B(n2583), 
	.A(\addr_calc/iir_read_calc/count[9] ));
   NAND4X1TS U3394 (.Y(n2784), 
	.D(n817), 
	.C(n816), 
	.B(n815), 
	.A(n814));
   NAND4X2TS U3395 (.Y(n2788), 
	.D(n918), 
	.C(n917), 
	.B(n916), 
	.A(n915));
   NOR4XLTS U3396 (.Y(n916), 
	.D(n2039), 
	.C(\addr_calc/iir_write_calc/count[7] ), 
	.B(n2041), 
	.A(n2562));
   NAND4X1TS U3397 (.Y(n2789), 
	.D(n922), 
	.C(n921), 
	.B(n920), 
	.A(n919));
endmodule

