library verilog;
use verilog.vl_types.all;
entity addr_calc_top_tb is
end addr_calc_top_tb;
