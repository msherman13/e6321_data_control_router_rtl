library verilog;
use verilog.vl_types.all;
entity dc_router_top_tb is
end dc_router_top_tb;
