library verilog;
use verilog.vl_types.all;
entity fft_addr_calc_tb is
end fft_addr_calc_tb;
