
module counter1 ( filesize, enable, pause, clk, count, done );
  input [31:0] filesize;
  output [31:0] count;
  input enable, pause, clk;
  output done;
  wire   N38, N43, N44, N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55,
         N56, N57, N58, N59, N60, N61, N62, N63, N64, N65, N66, N67, N68, N69,
         N70, N71, N72, N73, N74, n4, n5, n6, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, \add_x_22_0/carry[2] ,
         \add_x_22_0/carry[3] , \add_x_22_0/carry[4] , \add_x_22_0/carry[5] ,
         \add_x_22_0/carry[6] , \add_x_22_0/carry[7] , \add_x_22_0/carry[8] ,
         \add_x_22_0/carry[9] , \add_x_22_0/carry[10] , \add_x_22_0/carry[11] ,
         \add_x_22_0/carry[12] , \add_x_22_0/carry[13] ,
         \add_x_22_0/carry[14] , \add_x_22_0/carry[15] ,
         \add_x_22_0/carry[16] , \add_x_22_0/carry[17] ,
         \add_x_22_0/carry[18] , \add_x_22_0/carry[19] ,
         \add_x_22_0/carry[20] , \add_x_22_0/carry[21] ,
         \add_x_22_0/carry[22] , \add_x_22_0/carry[23] ,
         \add_x_22_0/carry[24] , \add_x_22_0/carry[25] ,
         \add_x_22_0/carry[26] , \add_x_22_0/carry[27] ,
         \add_x_22_0/carry[28] , \add_x_22_0/carry[29] ,
         \add_x_22_0/carry[30] , \add_x_22_0/carry[31] , n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243;

  NAND4X1TS U41 ( .A(n12), .B(n13), .C(n14), .D(n15), .Y(n11) );
  NOR4XLTS U42 ( .A(count[30]), .B(count[2]), .C(count[29]), .D(count[28]), 
        .Y(n15) );
  NOR4XLTS U43 ( .A(count[27]), .B(count[26]), .C(count[25]), .D(count[24]), 
        .Y(n14) );
  NOR4XLTS U44 ( .A(count[9]), .B(count[8]), .C(count[7]), .D(count[6]), .Y(
        n13) );
  NOR4XLTS U45 ( .A(count[5]), .B(count[4]), .C(count[3]), .D(count[31]), .Y(
        n12) );
  NAND4X1TS U46 ( .A(n16), .B(n17), .C(n18), .D(n19), .Y(n10) );
  NOR4XLTS U47 ( .A(count[16]), .B(count[15]), .C(count[14]), .D(count[13]), 
        .Y(n19) );
  NOR4XLTS U48 ( .A(count[12]), .B(count[11]), .C(count[10]), .D(n161), .Y(n18) );
  NOR4XLTS U49 ( .A(count[23]), .B(count[22]), .C(count[21]), .D(count[20]), 
        .Y(n17) );
  NOR4XLTS U50 ( .A(count[1]), .B(count[19]), .C(count[18]), .D(count[17]), 
        .Y(n16) );
  DFFQX1TS \count_reg[31]  ( .D(n50), .CK(clk), .Q(count[31]) );
  DFFQX1TS \count_reg[29]  ( .D(n21), .CK(clk), .Q(count[29]) );
  DFFQX1TS \count_reg[26]  ( .D(n24), .CK(clk), .Q(count[26]) );
  DFFQX1TS \count_reg[30]  ( .D(n20), .CK(clk), .Q(count[30]) );
  DFFQX1TS \count_reg[25]  ( .D(n25), .CK(clk), .Q(count[25]) );
  DFFQX1TS \count_reg[22]  ( .D(n28), .CK(clk), .Q(count[22]) );
  DFFQX1TS \count_reg[20]  ( .D(n30), .CK(clk), .Q(count[20]) );
  DFFQX1TS \count_reg[24]  ( .D(n26), .CK(clk), .Q(count[24]) );
  DFFQX1TS \count_reg[28]  ( .D(n22), .CK(clk), .Q(count[28]) );
  DFFQX1TS \count_reg[16]  ( .D(n34), .CK(clk), .Q(count[16]) );
  DFFQX1TS \count_reg[23]  ( .D(n27), .CK(clk), .Q(count[23]) );
  DFFQX1TS \count_reg[27]  ( .D(n23), .CK(clk), .Q(count[27]) );
  DFFQX1TS \count_reg[14]  ( .D(n36), .CK(clk), .Q(count[14]) );
  DFFQX1TS \count_reg[18]  ( .D(n32), .CK(clk), .Q(count[18]) );
  DFFQX1TS \count_reg[21]  ( .D(n29), .CK(clk), .Q(count[21]) );
  DFFQX1TS \count_reg[8]  ( .D(n42), .CK(clk), .Q(count[8]) );
  DFFQX1TS \count_reg[11]  ( .D(n39), .CK(clk), .Q(count[11]) );
  DFFQX1TS \count_reg[15]  ( .D(n35), .CK(clk), .Q(count[15]) );
  DFFQX1TS \count_reg[19]  ( .D(n31), .CK(clk), .Q(count[19]) );
  DFFQX1TS \count_reg[17]  ( .D(n33), .CK(clk), .Q(count[17]) );
  DFFQX1TS \count_reg[7]  ( .D(n43), .CK(clk), .Q(count[7]) );
  DFFQX1TS \count_reg[10]  ( .D(n40), .CK(clk), .Q(count[10]) );
  DFFQX1TS \count_reg[4]  ( .D(n46), .CK(clk), .Q(count[4]) );
  DFFQX1TS \count_reg[6]  ( .D(n44), .CK(clk), .Q(count[6]) );
  DFFQX1TS \count_reg[13]  ( .D(n37), .CK(clk), .Q(count[13]) );
  DFFQX1TS \count_reg[5]  ( .D(n45), .CK(clk), .Q(count[5]) );
  DFFQX1TS \count_reg[9]  ( .D(n41), .CK(clk), .Q(count[9]) );
  DFFQX1TS \count_reg[12]  ( .D(n38), .CK(clk), .Q(count[12]) );
  DFFQX1TS \count_reg[3]  ( .D(n47), .CK(clk), .Q(count[3]) );
  DFFQX1TS \count_reg[2]  ( .D(n48), .CK(clk), .Q(count[2]) );
  DFFQX1TS \count_reg[1]  ( .D(n49), .CK(clk), .Q(count[1]) );
  NOR2X1TS U40 ( .A(n10), .B(n11), .Y(n6) );
  AOI21X1TS U38 ( .A0(n9), .A1(N38), .B0(n129), .Y(n4) );
  NOR3X1TS U35 ( .A(n234), .B(n6), .C(n129), .Y(n5) );
  ADDHXLTS \add_x_22_0/U1_1_30  ( .A(count[30]), .B(\add_x_22_0/carry[30] ), 
        .CO(\add_x_22_0/carry[31] ), .S(N73) );
  ADDHXLTS \add_x_22_0/U1_1_29  ( .A(count[29]), .B(\add_x_22_0/carry[29] ), 
        .CO(\add_x_22_0/carry[30] ), .S(N72) );
  ADDHXLTS \add_x_22_0/U1_1_28  ( .A(count[28]), .B(\add_x_22_0/carry[28] ), 
        .CO(\add_x_22_0/carry[29] ), .S(N71) );
  ADDHXLTS \add_x_22_0/U1_1_27  ( .A(count[27]), .B(\add_x_22_0/carry[27] ), 
        .CO(\add_x_22_0/carry[28] ), .S(N70) );
  ADDHXLTS \add_x_22_0/U1_1_26  ( .A(count[26]), .B(\add_x_22_0/carry[26] ), 
        .CO(\add_x_22_0/carry[27] ), .S(N69) );
  ADDHXLTS \add_x_22_0/U1_1_25  ( .A(count[25]), .B(\add_x_22_0/carry[25] ), 
        .CO(\add_x_22_0/carry[26] ), .S(N68) );
  ADDHXLTS \add_x_22_0/U1_1_24  ( .A(count[24]), .B(\add_x_22_0/carry[24] ), 
        .CO(\add_x_22_0/carry[25] ), .S(N67) );
  ADDHXLTS \add_x_22_0/U1_1_23  ( .A(count[23]), .B(\add_x_22_0/carry[23] ), 
        .CO(\add_x_22_0/carry[24] ), .S(N66) );
  ADDHXLTS \add_x_22_0/U1_1_22  ( .A(count[22]), .B(\add_x_22_0/carry[22] ), 
        .CO(\add_x_22_0/carry[23] ), .S(N65) );
  ADDHXLTS \add_x_22_0/U1_1_21  ( .A(count[21]), .B(\add_x_22_0/carry[21] ), 
        .CO(\add_x_22_0/carry[22] ), .S(N64) );
  ADDHXLTS \add_x_22_0/U1_1_20  ( .A(count[20]), .B(\add_x_22_0/carry[20] ), 
        .CO(\add_x_22_0/carry[21] ), .S(N63) );
  ADDHXLTS \add_x_22_0/U1_1_19  ( .A(count[19]), .B(\add_x_22_0/carry[19] ), 
        .CO(\add_x_22_0/carry[20] ), .S(N62) );
  ADDHXLTS \add_x_22_0/U1_1_18  ( .A(count[18]), .B(\add_x_22_0/carry[18] ), 
        .CO(\add_x_22_0/carry[19] ), .S(N61) );
  ADDHXLTS \add_x_22_0/U1_1_17  ( .A(count[17]), .B(\add_x_22_0/carry[17] ), 
        .CO(\add_x_22_0/carry[18] ), .S(N60) );
  ADDHXLTS \add_x_22_0/U1_1_16  ( .A(count[16]), .B(\add_x_22_0/carry[16] ), 
        .CO(\add_x_22_0/carry[17] ), .S(N59) );
  ADDHXLTS \add_x_22_0/U1_1_15  ( .A(count[15]), .B(\add_x_22_0/carry[15] ), 
        .CO(\add_x_22_0/carry[16] ), .S(N58) );
  ADDHXLTS \add_x_22_0/U1_1_14  ( .A(count[14]), .B(\add_x_22_0/carry[14] ), 
        .CO(\add_x_22_0/carry[15] ), .S(N57) );
  ADDHXLTS \add_x_22_0/U1_1_13  ( .A(count[13]), .B(\add_x_22_0/carry[13] ), 
        .CO(\add_x_22_0/carry[14] ), .S(N56) );
  ADDHXLTS \add_x_22_0/U1_1_12  ( .A(count[12]), .B(\add_x_22_0/carry[12] ), 
        .CO(\add_x_22_0/carry[13] ), .S(N55) );
  ADDHXLTS \add_x_22_0/U1_1_11  ( .A(count[11]), .B(\add_x_22_0/carry[11] ), 
        .CO(\add_x_22_0/carry[12] ), .S(N54) );
  ADDHXLTS \add_x_22_0/U1_1_10  ( .A(count[10]), .B(\add_x_22_0/carry[10] ), 
        .CO(\add_x_22_0/carry[11] ), .S(N53) );
  ADDHXLTS \add_x_22_0/U1_1_9  ( .A(count[9]), .B(\add_x_22_0/carry[9] ), .CO(
        \add_x_22_0/carry[10] ), .S(N52) );
  ADDHXLTS \add_x_22_0/U1_1_8  ( .A(count[8]), .B(\add_x_22_0/carry[8] ), .CO(
        \add_x_22_0/carry[9] ), .S(N51) );
  ADDHXLTS \add_x_22_0/U1_1_7  ( .A(count[7]), .B(\add_x_22_0/carry[7] ), .CO(
        \add_x_22_0/carry[8] ), .S(N50) );
  ADDHXLTS \add_x_22_0/U1_1_6  ( .A(count[6]), .B(\add_x_22_0/carry[6] ), .CO(
        \add_x_22_0/carry[7] ), .S(N49) );
  ADDHXLTS \add_x_22_0/U1_1_5  ( .A(count[5]), .B(\add_x_22_0/carry[5] ), .CO(
        \add_x_22_0/carry[6] ), .S(N48) );
  ADDHXLTS \add_x_22_0/U1_1_4  ( .A(count[4]), .B(\add_x_22_0/carry[4] ), .CO(
        \add_x_22_0/carry[5] ), .S(N47) );
  ADDHXLTS \add_x_22_0/U1_1_3  ( .A(count[3]), .B(\add_x_22_0/carry[3] ), .CO(
        \add_x_22_0/carry[4] ), .S(N46) );
  ADDHXLTS \add_x_22_0/U1_1_2  ( .A(count[2]), .B(\add_x_22_0/carry[2] ), .CO(
        \add_x_22_0/carry[3] ), .S(N45) );
  ADDHXLTS \add_x_22_0/U1_1_1  ( .A(count[1]), .B(count[0]), .CO(
        \add_x_22_0/carry[2] ), .S(N44) );
  AO22XLTS U22 ( .A0(n238), .A1(count[12]), .B0(n5), .B1(N55), .Y(n38) );
  AO22XLTS U4 ( .A0(n4), .A1(count[30]), .B0(n233), .B1(N73), .Y(n20) );
  AO22XLTS U6 ( .A0(n234), .A1(count[28]), .B0(n231), .B1(N71), .Y(n22) );
  AO22XLTS U20 ( .A0(n241), .A1(count[14]), .B0(n232), .B1(N57), .Y(n36) );
  AO22XLTS U19 ( .A0(n4), .A1(count[15]), .B0(n232), .B1(N58), .Y(n35) );
  AO22XLTS U21 ( .A0(n243), .A1(count[13]), .B0(n232), .B1(N56), .Y(n37) );
  AO22XLTS U5 ( .A0(n234), .A1(count[29]), .B0(n233), .B1(N72), .Y(n21) );
  AO22XLTS U34 ( .A0(n240), .A1(count[31]), .B0(n225), .B1(N74), .Y(n50) );
  AO22XLTS U16 ( .A0(n237), .A1(count[18]), .B0(n228), .B1(N61), .Y(n32) );
  AO22XLTS U33 ( .A0(n243), .A1(count[1]), .B0(n225), .B1(N44), .Y(n49) );
  AO22XLTS U32 ( .A0(n240), .A1(count[2]), .B0(n225), .B1(N45), .Y(n48) );
  AO22XLTS U7 ( .A0(n235), .A1(count[27]), .B0(n230), .B1(N70), .Y(n23) );
  AO22XLTS U8 ( .A0(n235), .A1(count[26]), .B0(n230), .B1(N69), .Y(n24) );
  AO22XLTS U31 ( .A0(n240), .A1(count[3]), .B0(n225), .B1(N46), .Y(n47) );
  AO22XLTS U9 ( .A0(n235), .A1(count[25]), .B0(n230), .B1(N68), .Y(n25) );
  AO22XLTS U10 ( .A0(n235), .A1(count[24]), .B0(n230), .B1(N67), .Y(n26) );
  AO22XLTS U30 ( .A0(n243), .A1(count[4]), .B0(n226), .B1(N47), .Y(n46) );
  AO22XLTS U11 ( .A0(n236), .A1(count[23]), .B0(n229), .B1(N66), .Y(n27) );
  AO22XLTS U12 ( .A0(n236), .A1(count[22]), .B0(n229), .B1(N65), .Y(n28) );
  AO22XLTS U29 ( .A0(n239), .A1(count[5]), .B0(n226), .B1(N48), .Y(n45) );
  AO22XLTS U13 ( .A0(n236), .A1(count[21]), .B0(n229), .B1(N64), .Y(n29) );
  AO22XLTS U14 ( .A0(n236), .A1(count[20]), .B0(n229), .B1(N63), .Y(n30) );
  AO22XLTS U28 ( .A0(n239), .A1(count[6]), .B0(n226), .B1(N49), .Y(n44) );
  AO22XLTS U24 ( .A0(n238), .A1(count[10]), .B0(n227), .B1(N53), .Y(n40) );
  AO22XLTS U27 ( .A0(n239), .A1(count[7]), .B0(n226), .B1(N50), .Y(n43) );
  AO22XLTS U18 ( .A0(n237), .A1(count[16]), .B0(n228), .B1(N59), .Y(n34) );
  AO22XLTS U15 ( .A0(n237), .A1(count[19]), .B0(n228), .B1(N62), .Y(n31) );
  AO22XLTS U26 ( .A0(n239), .A1(count[8]), .B0(n227), .B1(N51), .Y(n42) );
  AO22XLTS U17 ( .A0(n237), .A1(count[17]), .B0(n228), .B1(N60), .Y(n33) );
  AO22XLTS U23 ( .A0(n238), .A1(count[11]), .B0(n227), .B1(N54), .Y(n39) );
  AO22XLTS U25 ( .A0(n238), .A1(count[9]), .B0(n227), .B1(N52), .Y(n41) );
  SDFFXLTS done_reg ( .D(N38), .SI(1'b1), .SE(n129), .CK(clk), .QN(done) );
  DFFXLTS \count_reg[0]  ( .D(n51), .CK(clk), .Q(count[0]), .QN(N43) );
  NOR4XLTS U52 ( .A(n137), .B(n139), .C(n157), .D(n159), .Y(n191) );
  XNOR2X1TS U53 ( .A(n104), .B(count[17]), .Y(n52) );
  XOR2X1TS U54 ( .A(n122), .B(count[19]), .Y(n53) );
  XOR2X1TS U55 ( .A(n149), .B(count[18]), .Y(n54) );
  OAI211X1TS U56 ( .A0(n53), .A1(n149), .B0(n203), .C0(n54), .Y(n55) );
  AO21X1TS U57 ( .A0(n53), .A1(n149), .B0(n55), .Y(n56) );
  OAI31X1TS U58 ( .A0(n53), .A1(n203), .A2(n54), .B0(n56), .Y(n57) );
  XOR2X1TS U59 ( .A(n108), .B(count[11]), .Y(n58) );
  XOR2X1TS U60 ( .A(n120), .B(count[15]), .Y(n59) );
  XOR2X1TS U61 ( .A(n145), .B(count[14]), .Y(n60) );
  OAI211X1TS U62 ( .A0(n59), .A1(n145), .B0(n183), .C0(n60), .Y(n61) );
  AO21X1TS U63 ( .A0(n59), .A1(n145), .B0(n61), .Y(n62) );
  OAI31X1TS U64 ( .A0(n59), .A1(n183), .A2(n60), .B0(n62), .Y(n63) );
  XOR2X1TS U65 ( .A(n112), .B(count[8]), .Y(n64) );
  XOR2X1TS U66 ( .A(n124), .B(count[13]), .Y(n65) );
  XOR2X1TS U67 ( .A(n147), .B(count[12]), .Y(n66) );
  OAI211X1TS U68 ( .A0(n65), .A1(n147), .B0(n184), .C0(n66), .Y(n67) );
  AO21X1TS U69 ( .A0(n65), .A1(n147), .B0(n67), .Y(n68) );
  OAI31X1TS U70 ( .A0(n65), .A1(n184), .A2(n66), .B0(n68), .Y(n69) );
  XOR2X1TS U71 ( .A(n116), .B(count[5]), .Y(n70) );
  XOR2X1TS U72 ( .A(n128), .B(count[10]), .Y(n71) );
  XOR2X1TS U73 ( .A(n141), .B(count[9]), .Y(n72) );
  OAI211X1TS U74 ( .A0(n71), .A1(n141), .B0(n185), .C0(n72), .Y(n73) );
  AO21X1TS U75 ( .A0(n71), .A1(n141), .B0(n73), .Y(n74) );
  OAI31X1TS U76 ( .A0(n71), .A1(n185), .A2(n72), .B0(n74), .Y(n75) );
  XNOR2X1TS U77 ( .A(count[2]), .B(n139), .Y(n76) );
  NOR2X1TS U78 ( .A(n157), .B(n160), .Y(n77) );
  OAI31X1TS U79 ( .A0(n190), .A1(n188), .A2(n189), .B0(n187), .Y(n78) );
  OAI21X1TS U80 ( .A0(n76), .A1(n77), .B0(n78), .Y(n79) );
  AOI211X1TS U81 ( .A0(n76), .A1(n77), .B0(n199), .C0(n79), .Y(n80) );
  OAI211X1TS U82 ( .A0(n200), .A1(n70), .B0(n80), .C0(n75), .Y(n81) );
  AOI21X1TS U83 ( .A0(n200), .A1(n70), .B0(n81), .Y(n82) );
  OAI211X1TS U84 ( .A0(n201), .A1(n64), .B0(n82), .C0(n69), .Y(n83) );
  AOI21X1TS U85 ( .A0(n201), .A1(n64), .B0(n83), .Y(n84) );
  OAI211X1TS U86 ( .A0(n202), .A1(n58), .B0(n84), .C0(n63), .Y(n85) );
  AOI21X1TS U87 ( .A0(n202), .A1(n58), .B0(n85), .Y(n86) );
  OAI211X1TS U88 ( .A0(n52), .A1(n204), .B0(n86), .C0(n57), .Y(n87) );
  AOI21X1TS U89 ( .A0(n52), .A1(n204), .B0(n87), .Y(n88) );
  XNOR2X1TS U90 ( .A(n182), .B(count[16]), .Y(n89) );
  NAND2X1TS U91 ( .A(n135), .B(n89), .Y(n90) );
  OAI211X1TS U92 ( .A0(n135), .A1(n89), .B0(n88), .C0(n90), .Y(n205) );
  CLKINVX1TS U93 ( .A(n234), .Y(n91) );
  OAI21X1TS U94 ( .A0(n6), .A1(N43), .B0(n91), .Y(n92) );
  OAI2BB2XLTS U95 ( .B0(n129), .B1(n92), .A0N(n240), .A1N(n161), .Y(n51) );
  OAI211XLTS U97 ( .A0(n219), .A1(n218), .B0(n217), .C0(n216), .Y(n220) );
  OAI211XLTS U98 ( .A0(n214), .A1(n213), .B0(n212), .C0(n211), .Y(n215) );
  OAI31XLTS U99 ( .A0(n171), .A1(n170), .A2(n169), .B0(n168), .Y(n217) );
  OAI211XLTS U100 ( .A0(n209), .A1(n208), .B0(n207), .C0(n206), .Y(n210) );
  AOI21XLTS U101 ( .A0(n209), .A1(n208), .B0(n205), .Y(n206) );
  OAI31XLTS U102 ( .A0(n176), .A1(n175), .A2(n174), .B0(n173), .Y(n212) );
  OAI211XLTS U103 ( .A0(n171), .A1(n143), .B0(n170), .C0(n169), .Y(n167) );
  OAI211XLTS U104 ( .A0(n176), .A1(n155), .B0(n175), .C0(n174), .Y(n172) );
  AOI221XLTS U105 ( .A0(n195), .A1(n133), .B0(n194), .B1(n137), .C0(n193), .Y(
        n198) );
  OAI22XLTS U106 ( .A0(n133), .A1(n195), .B0(n194), .B1(n137), .Y(n193) );
  MXI2XLTS U107 ( .A(count[0]), .B(n159), .S0(n196), .Y(n197) );
  XOR2XLTS U108 ( .A(n151), .B(count[6]), .Y(n189) );
  NOR3XLTS U109 ( .A(n139), .B(n157), .C(n160), .Y(n192) );
  XOR2XLTS U110 ( .A(n157), .B(count[1]), .Y(n196) );
  INVX1TS U111 ( .A(n158), .Y(n159) );
  INVX1TS U112 ( .A(n99), .Y(n100) );
  INVX1TS U113 ( .A(n115), .Y(n116) );
  INVX1TS U114 ( .A(n127), .Y(n128) );
  INVX1TS U115 ( .A(n123), .Y(n124) );
  INVX1TS U116 ( .A(n146), .Y(n147) );
  INVX1TS U117 ( .A(n119), .Y(n120) );
  INVX1TS U118 ( .A(n136), .Y(n137) );
  INVX1TS U119 ( .A(n132), .Y(n133) );
  INVX1TS U120 ( .A(n138), .Y(n139) );
  INVX1TS U121 ( .A(n144), .Y(n145) );
  INVX1TS U122 ( .A(n134), .Y(n135) );
  INVX2TS U123 ( .A(n156), .Y(n157) );
  INVX1TS U124 ( .A(n103), .Y(n104) );
  INVX1TS U125 ( .A(n111), .Y(n112) );
  INVX1TS U126 ( .A(n121), .Y(n122) );
  INVX2TS U127 ( .A(n148), .Y(n149) );
  INVX2TS U128 ( .A(n150), .Y(n151) );
  INVX2TS U129 ( .A(n152), .Y(n153) );
  INVX2TS U130 ( .A(n154), .Y(n155) );
  CLKINVX2TS U131 ( .A(n125), .Y(n126) );
  CLKINVX2TS U132 ( .A(n130), .Y(n131) );
  CLKINVX2TS U133 ( .A(n117), .Y(n118) );
  INVX2TS U134 ( .A(n142), .Y(n143) );
  INVX1TS U135 ( .A(n113), .Y(n114) );
  INVX1TS U136 ( .A(n95), .Y(n96) );
  INVX1TS U137 ( .A(n101), .Y(n102) );
  INVX1TS U138 ( .A(n109), .Y(n110) );
  INVX1TS U139 ( .A(n105), .Y(n106) );
  INVX1TS U140 ( .A(n97), .Y(n98) );
  INVX1TS U141 ( .A(n140), .Y(n141) );
  INVX1TS U142 ( .A(n107), .Y(n108) );
  INVXLTS U143 ( .A(filesize[31]), .Y(n95) );
  INVXLTS U144 ( .A(pause), .Y(n9) );
  INVXLTS U145 ( .A(filesize[21]), .Y(n97) );
  INVXLTS U146 ( .A(filesize[7]), .Y(n99) );
  INVXLTS U147 ( .A(filesize[25]), .Y(n101) );
  INVXLTS U148 ( .A(filesize[17]), .Y(n103) );
  INVXLTS U149 ( .A(filesize[22]), .Y(n105) );
  INVXLTS U150 ( .A(filesize[11]), .Y(n107) );
  INVXLTS U151 ( .A(filesize[23]), .Y(n109) );
  INVXLTS U152 ( .A(filesize[8]), .Y(n111) );
  INVXLTS U153 ( .A(filesize[26]), .Y(n113) );
  INVXLTS U154 ( .A(filesize[5]), .Y(n115) );
  INVXLTS U155 ( .A(filesize[29]), .Y(n117) );
  INVXLTS U156 ( .A(filesize[15]), .Y(n119) );
  INVXLTS U157 ( .A(filesize[19]), .Y(n121) );
  INVXLTS U158 ( .A(filesize[13]), .Y(n123) );
  INVXLTS U159 ( .A(filesize[28]), .Y(n125) );
  INVXLTS U160 ( .A(filesize[10]), .Y(n127) );
  INVXLTS U161 ( .A(enable), .Y(n129) );
  INVXLTS U162 ( .A(filesize[30]), .Y(n130) );
  INVXLTS U163 ( .A(filesize[4]), .Y(n132) );
  INVXLTS U164 ( .A(filesize[16]), .Y(n134) );
  INVXLTS U165 ( .A(filesize[3]), .Y(n136) );
  INVXLTS U166 ( .A(filesize[2]), .Y(n138) );
  INVXLTS U167 ( .A(filesize[9]), .Y(n140) );
  INVXLTS U168 ( .A(filesize[27]), .Y(n142) );
  INVXLTS U169 ( .A(filesize[14]), .Y(n144) );
  INVXLTS U170 ( .A(filesize[12]), .Y(n146) );
  INVXLTS U171 ( .A(filesize[18]), .Y(n148) );
  INVXLTS U172 ( .A(filesize[6]), .Y(n150) );
  INVXLTS U173 ( .A(filesize[20]), .Y(n152) );
  INVXLTS U174 ( .A(filesize[24]), .Y(n154) );
  INVXLTS U175 ( .A(filesize[1]), .Y(n156) );
  INVXLTS U176 ( .A(filesize[0]), .Y(n158) );
  INVXLTS U177 ( .A(n158), .Y(n160) );
  INVX2TS U178 ( .A(N43), .Y(n161) );
  OAI211XLTS U179 ( .A0(count[0]), .A1(n159), .B0(n198), .C0(n197), .Y(n199)
         );
  XOR2X1TS U180 ( .A(\add_x_22_0/carry[31] ), .B(count[31]), .Y(N74) );
  XOR2X1TS U181 ( .A(n96), .B(count[31]), .Y(n166) );
  XOR2X1TS U182 ( .A(n131), .B(count[30]), .Y(n165) );
  XOR2X1TS U183 ( .A(n114), .B(count[26]), .Y(n218) );
  XOR2X1TS U184 ( .A(n126), .B(count[28]), .Y(n171) );
  XOR2X1TS U185 ( .A(n143), .B(count[27]), .Y(n170) );
  AO21X1TS U186 ( .A0(n171), .A1(n143), .B0(n167), .Y(n168) );
  XOR2X1TS U187 ( .A(n110), .B(count[23]), .Y(n213) );
  XOR2X1TS U188 ( .A(n102), .B(count[25]), .Y(n176) );
  XOR2X1TS U189 ( .A(n155), .B(count[24]), .Y(n175) );
  AO21X1TS U190 ( .A0(n176), .A1(n155), .B0(n172), .Y(n173) );
  XOR2X1TS U191 ( .A(n106), .B(count[22]), .Y(n208) );
  XOR2X1TS U192 ( .A(n98), .B(count[21]), .Y(n181) );
  XOR2X1TS U193 ( .A(n153), .B(count[20]), .Y(n180) );
  AO21X1TS U194 ( .A0(n181), .A1(n153), .B0(n177), .Y(n178) );
  XOR2X1TS U195 ( .A(n100), .B(count[7]), .Y(n190) );
  AO21X1TS U196 ( .A0(n190), .A1(n151), .B0(n186), .Y(n187) );
  XNOR2X1TS U197 ( .A(n191), .B(count[4]), .Y(n195) );
  XNOR2X1TS U198 ( .A(n192), .B(count[3]), .Y(n194) );
  XOR2X1TS U199 ( .A(n118), .B(count[29]), .Y(n223) );
  NOR2X1TS U200 ( .A(n118), .B(n224), .Y(n164) );
  OAI211X1TS U201 ( .A0(n166), .A1(n131), .B0(n165), .C0(n164), .Y(n162) );
  OAI31X1TS U202 ( .A0(n166), .A1(n165), .A2(n164), .B0(n163), .Y(n222) );
  AOI21X1TS U203 ( .A0(n219), .A1(n218), .B0(n215), .Y(n216) );
  AOI21X1TS U204 ( .A0(n224), .A1(n223), .B0(n220), .Y(n221) );
  OAI211X1TS U205 ( .A0(n224), .A1(n223), .B0(n222), .C0(n221), .Y(N38) );
  AOI21X1TS U206 ( .A0(n214), .A1(n213), .B0(n210), .Y(n211) );
  AO21X1TS U207 ( .A0(n166), .A1(n131), .B0(n162), .Y(n163) );
  NAND2BX1TS U208 ( .AN(n133), .B(n191), .Y(n200) );
  NOR3BX1TS U209 ( .AN(n183), .B(n120), .C(n145), .Y(n182) );
  NOR2BX1TS U210 ( .AN(n182), .B(n135), .Y(n204) );
  NOR2BX1TS U211 ( .AN(n204), .B(n104), .Y(n203) );
  OR2X2TS U212 ( .A(n106), .B(n209), .Y(n214) );
  NAND3BX1TS U213 ( .AN(n143), .B(n169), .C(n125), .Y(n224) );
  NOR2X1TS U214 ( .A(n108), .B(n202), .Y(n184) );
  NOR3BX1TS U215 ( .AN(n184), .B(n124), .C(n147), .Y(n183) );
  NAND3BX1TS U216 ( .AN(n98), .B(n179), .C(n152), .Y(n209) );
  NAND3BX1TS U217 ( .AN(n102), .B(n174), .C(n154), .Y(n219) );
  NOR2X1TS U218 ( .A(n114), .B(n219), .Y(n169) );
  NOR2X1TS U219 ( .A(n116), .B(n200), .Y(n188) );
  NAND3BX1TS U220 ( .AN(n100), .B(n188), .C(n150), .Y(n201) );
  NOR2X1TS U221 ( .A(n112), .B(n201), .Y(n185) );
  NAND3BX1TS U222 ( .AN(n141), .B(n185), .C(n127), .Y(n202) );
  NOR3BX1TS U223 ( .AN(n203), .B(n122), .C(n149), .Y(n179) );
  NOR2X1TS U224 ( .A(n110), .B(n214), .Y(n174) );
  OAI211XLTS U225 ( .A0(n181), .A1(n153), .B0(n180), .C0(n179), .Y(n177) );
  OAI31XLTS U226 ( .A0(n181), .A1(n180), .A2(n179), .B0(n178), .Y(n207) );
  OAI211XLTS U227 ( .A0(n190), .A1(n151), .B0(n189), .C0(n188), .Y(n186) );
  CLKBUFX2TS U228 ( .A(n243), .Y(n234) );
  CLKBUFX2TS U229 ( .A(n4), .Y(n243) );
  CLKBUFX2TS U230 ( .A(n242), .Y(n241) );
  CLKBUFX2TS U231 ( .A(n4), .Y(n242) );
  CLKBUFX2TS U232 ( .A(n5), .Y(n233) );
  CLKBUFX2TS U233 ( .A(n232), .Y(n227) );
  CLKBUFX2TS U234 ( .A(n241), .Y(n238) );
  CLKBUFX2TS U235 ( .A(n233), .Y(n225) );
  CLKBUFX2TS U236 ( .A(n241), .Y(n239) );
  CLKBUFX2TS U237 ( .A(n233), .Y(n226) );
  CLKBUFX2TS U238 ( .A(n231), .Y(n228) );
  CLKBUFX2TS U239 ( .A(n241), .Y(n237) );
  CLKBUFX2TS U240 ( .A(n231), .Y(n229) );
  CLKBUFX2TS U241 ( .A(n242), .Y(n236) );
  CLKBUFX2TS U242 ( .A(n242), .Y(n235) );
  CLKBUFX2TS U243 ( .A(n5), .Y(n231) );
  CLKBUFX2TS U244 ( .A(n5), .Y(n232) );
  CLKBUFX2TS U245 ( .A(n231), .Y(n230) );
  CLKBUFX2TS U246 ( .A(n242), .Y(n240) );
endmodule

