library verilog;
use verilog.vl_types.all;
entity pla_top_tb is
end pla_top_tb;
