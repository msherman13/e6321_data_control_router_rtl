library verilog;
use verilog.vl_types.all;
entity data_bus_controller_tb is
end data_bus_controller_tb;
